* ---- BEGIN sky130_fd_pr__nfet_01v8__subvt_mismatch.corner.spice ----
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8__toxe_slope=3.443e-03
.param sky130_fd_pr__nfet_01v8__lint_slope=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_slope=0.11
.param sky130_fd_pr__nfet_01v8__voff_slope=0.015
.param sky130_fd_pr__nfet_01v8__vth0_slope=8.556e-03
.param sky130_fd_pr__nfet_01v8__vth0_slope1=1.0056e-02
.param sky130_fd_pr__nfet_01v8__wint_slope=0
* ---- END sky130_fd_pr__nfet_01v8__subvt_mismatch.corner.spice ----

* ---- BEGIN sky130_fd_pr__pfet_01v8__subvt_mismatch.corner.spice ----
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8__toxe_slope=4.443e-03
.param sky130_fd_pr__pfet_01v8__toxe_slope1=6.443e-03
.param sky130_fd_pr__pfet_01v8__toxe_slope2=3.443e-03
.param sky130_fd_pr__pfet_01v8__lint_slope=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope=0.1
.param sky130_fd_pr__pfet_01v8__nfactor_slope1=0.1
.param sky130_fd_pr__pfet_01v8__nfactor_slope2=0.0
.param sky130_fd_pr__pfet_01v8__voff_slope=0.015
.param sky130_fd_pr__pfet_01v8__voff_slope1=0.015
.param sky130_fd_pr__pfet_01v8__voff_slope2=0.017
.param sky130_fd_pr__pfet_01v8__vth0_slope=8.856e-03
.param sky130_fd_pr__pfet_01v8__vth0_slope1=1.0356e-02
.param sky130_fd_pr__pfet_01v8__vth0_slope2=7.356e-03
.param sky130_fd_pr__pfet_01v8__wint_slope=0

* ---- END sky130_fd_pr__pfet_01v8__subvt_mismatch.corner.spice ----

* ============================================================
* === ROOTCAUSE_UI_BEGIN ===
* ROOT-CAUSE OVERRIDES (USER / UI CONTROL)
* ============================================================
.param MC_MM_SWITCH = 1

.param X_cd     = 0
.param X_damage = 0
.param X_eot    = 0
.param X_act    = 0
.param X_rc     = 0

.param a_dlc  = 1.0e-9
.param a_dwc  = 0.0
.param a_toxe = 0.010
.param a_vth  = 0.020
.param a_u0   = 5.0e-4
.param a_nf   = 0.020
.param a_voff = 0.010
.param a_rdsw = 100

.param NP_SPLIT = 0

.param a_dlc_n  = 1.0e-9
.param a_dwc_n  = 0.0
.param a_toxe_n = 0.010
.param a_vth_n  = 0.020
.param a_u0_n   = 5.0e-4
.param a_nf_n   = 0.020
.param a_voff_n = 0.010
.param a_rdsw_n = 100

.param a_dlc_p  = 1.0e-9
.param a_dwc_p  = 0.0
.param a_toxe_p = 0.010
.param a_vth_p  = 0.020
.param a_u0_p   = 5.0e-4
.param a_nf_p   = 0.020
.param a_voff_p = 0.010
.param a_rdsw_p = 100

* ngspice ternary: cond ? a : b
.param A_DLC_N  = {NP_SPLIT ? a_dlc_n  : a_dlc}
.param A_DWC_N  = {NP_SPLIT ? a_dwc_n  : a_dwc}
.param A_TOXE_N = {NP_SPLIT ? a_toxe_n : a_toxe}
.param A_VTH_N  = {NP_SPLIT ? a_vth_n  : a_vth}
.param A_U0_N   = {NP_SPLIT ? a_u0_n   : a_u0}
.param A_NF_N   = {NP_SPLIT ? a_nf_n   : a_nf}
.param A_VOFF_N = {NP_SPLIT ? a_voff_n : a_voff}
.param A_RDSW_N = {NP_SPLIT ? a_rdsw_n : a_rdsw}

.param A_DLC_P  = {NP_SPLIT ? a_dlc_p  : a_dlc}
.param A_DWC_P  = {NP_SPLIT ? a_dwc_p  : a_dwc}
.param A_TOXE_P = {NP_SPLIT ? a_toxe_p : a_toxe}
.param A_VTH_P  = {NP_SPLIT ? a_vth_p  : a_vth}
.param A_U0_P   = {NP_SPLIT ? a_u0_p   : a_u0}
.param A_NF_P   = {NP_SPLIT ? a_nf_p   : a_nf}
.param A_VOFF_P = {NP_SPLIT ? a_voff_p : a_voff}
.param A_RDSW_P = {NP_SPLIT ? a_rdsw_p : a_rdsw}

* GLOBAL knobs
.param sky130_fd_pr__nfet_01v8__dlc_diff = {sky130_fd_pr__nfet_01v8__dlc_diff + A_DLC_N*X_cd}
.param sky130_fd_pr__nfet_01v8__dwc_diff = {sky130_fd_pr__nfet_01v8__dwc_diff + A_DWC_N*X_cd}
.param sky130_fd_pr__pfet_01v8__dlc_diff = {sky130_fd_pr__pfet_01v8__dlc_diff + A_DLC_P*X_cd}
.param sky130_fd_pr__pfet_01v8__dwc_diff = {sky130_fd_pr__pfet_01v8__dwc_diff + A_DWC_P*X_cd}

.param sky130_fd_pr__nfet_01v8__toxe_mult = {sky130_fd_pr__nfet_01v8__toxe_mult*(1 + A_TOXE_N*X_eot)}
.param sky130_fd_pr__pfet_01v8__toxe_mult = {sky130_fd_pr__pfet_01v8__toxe_mult*(1 + A_TOXE_P*X_eot)}

* BIN indexed knobs (0..3 example)
.param sky130_fd_pr__nfet_01v8__vth0_diff_0 = {sky130_fd_pr__nfet_01v8__vth0_diff_0 + A_VTH_N*X_act}
.param sky130_fd_pr__pfet_01v8__vth0_diff_0 = {sky130_fd_pr__pfet_01v8__vth0_diff_0 + A_VTH_P*X_act}
.param sky130_fd_pr__nfet_01v8__vth0_diff_1 = {sky130_fd_pr__nfet_01v8__vth0_diff_1 + A_VTH_N*X_act}
.param sky130_fd_pr__pfet_01v8__vth0_diff_1 = {sky130_fd_pr__pfet_01v8__vth0_diff_1 + A_VTH_P*X_act}
.param sky130_fd_pr__nfet_01v8__vth0_diff_2 = {sky130_fd_pr__nfet_01v8__vth0_diff_2 + A_VTH_N*X_act}
.param sky130_fd_pr__pfet_01v8__vth0_diff_2 = {sky130_fd_pr__pfet_01v8__vth0_diff_2 + A_VTH_P*X_act}
.param sky130_fd_pr__nfet_01v8__vth0_diff_3 = {sky130_fd_pr__nfet_01v8__vth0_diff_3 + A_VTH_N*X_act}
.param sky130_fd_pr__pfet_01v8__vth0_diff_3 = {sky130_fd_pr__pfet_01v8__vth0_diff_3 + A_VTH_P*X_act}

.param sky130_fd_pr__nfet_01v8__u0_diff_0 = {sky130_fd_pr__nfet_01v8__u0_diff_0 - A_U0_N*X_damage}
.param sky130_fd_pr__pfet_01v8__u0_diff_0 = {sky130_fd_pr__pfet_01v8__u0_diff_0 - A_U0_P*X_damage}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_0 = {sky130_fd_pr__nfet_01v8__nfactor_diff_0 + A_NF_N*X_damage}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_0 = {sky130_fd_pr__pfet_01v8__nfactor_diff_0 + A_NF_P*X_damage}
.param sky130_fd_pr__nfet_01v8__voff_diff_0 = {sky130_fd_pr__nfet_01v8__voff_diff_0 + A_VOFF_N*X_damage}
.param sky130_fd_pr__pfet_01v8__voff_diff_0 = {sky130_fd_pr__pfet_01v8__voff_diff_0 + A_VOFF_P*X_damage}

.param sky130_fd_pr__nfet_01v8__rdsw_diff_0 = {sky130_fd_pr__nfet_01v8__rdsw_diff_0 + A_RDSW_N*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_0 = {sky130_fd_pr__pfet_01v8__rdsw_diff_0 + A_RDSW_P*X_rc}

* ============================================================
* END ROOT-CAUSE OVERRIDES
* === ROOTCAUSE_UI_END ===
* ============================================================
