* ---- BEGIN sky130_fd_pr__nfet_01v8__subvt_mismatch.corner.spice ----
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8__toxe_slope=3.443e-03
.param sky130_fd_pr__nfet_01v8__lint_slope=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_slope=0.11
.param sky130_fd_pr__nfet_01v8__voff_slope=0.015
.param sky130_fd_pr__nfet_01v8__vth0_slope=8.556e-03
.param sky130_fd_pr__nfet_01v8__vth0_slope1=1.0056e-02
.param sky130_fd_pr__nfet_01v8__wint_slope=0
* ---- END sky130_fd_pr__nfet_01v8__subvt_mismatch.corner.spice ----

* ---- BEGIN sky130_fd_pr__pfet_01v8__subvt_mismatch.corner.spice ----
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8__toxe_slope=4.443e-03
.param sky130_fd_pr__pfet_01v8__toxe_slope1=6.443e-03
.param sky130_fd_pr__pfet_01v8__toxe_slope2=3.443e-03
.param sky130_fd_pr__pfet_01v8__lint_slope=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope=0.1
.param sky130_fd_pr__pfet_01v8__nfactor_slope1=0.1
.param sky130_fd_pr__pfet_01v8__nfactor_slope2=0.0
.param sky130_fd_pr__pfet_01v8__voff_slope=0.015
.param sky130_fd_pr__pfet_01v8__voff_slope1=0.015
.param sky130_fd_pr__pfet_01v8__voff_slope2=0.017
.param sky130_fd_pr__pfet_01v8__vth0_slope=8.856e-03
.param sky130_fd_pr__pfet_01v8__vth0_slope1=1.0356e-02
.param sky130_fd_pr__pfet_01v8__vth0_slope2=7.356e-03
.param sky130_fd_pr__pfet_01v8__wint_slope=0

* ---- END sky130_fd_pr__pfet_01v8__subvt_mismatch.corner.spice ----

* ============================================================
* === ROOTCAUSE_UI_BEGIN ===
* ROOT-CAUSE OVERRIDES (USER / UI CONTROL)
* Auto-generated: full wafer variable mapping to latent X variables
* ============================================================
.param MC_MM_SWITCH = 1

.param X_cd     = 0
.param X_damage = 0
.param X_eot    = 0
.param X_act    = 0
.param X_rc     = 0

.param a_dlc  = 1.0e-9
.param a_dwc  = 0.0
.param a_toxe = 0.010
.param a_vth  = 0.020
.param a_u0   = 5.0e-4
.param a_nf   = 0.020
.param a_voff = 0.010
.param a_rdsw = 100

.param NP_SPLIT = 0

.param a_dlc_n = 1.0e-9
.param a_dwc_n = 0.0
.param a_toxe_n = 0.010
.param a_vth_n = 0.020
.param a_u0_n = 5.0e-4
.param a_nf_n = 0.020
.param a_voff_n = 0.010
.param a_rdsw_n = 100
.param a_dlc_p = 1.0e-9
.param a_dwc_p = 0.0
.param a_toxe_p = 0.010
.param a_vth_p = 0.020
.param a_u0_p = 5.0e-4
.param a_nf_p = 0.020
.param a_voff_p = 0.010
.param a_rdsw_p = 100

* Legacy UI aliases
.param A_DLC_N  = {NP_SPLIT ? a_dlc_n  : a_dlc}
.param A_DWC_N  = {NP_SPLIT ? a_dwc_n  : a_dwc}
.param A_TOXE_N = {NP_SPLIT ? a_toxe_n : a_toxe}
.param A_VTH_N  = {NP_SPLIT ? a_vth_n  : a_vth}
.param A_U0_N   = {NP_SPLIT ? a_u0_n   : a_u0}
.param A_NF_N   = {NP_SPLIT ? a_nf_n   : a_nf}
.param A_VOFF_N = {NP_SPLIT ? a_voff_n : a_voff}
.param A_RDSW_N = {NP_SPLIT ? a_rdsw_n : a_rdsw}
.param A_DLC_P  = {NP_SPLIT ? a_dlc_p  : a_dlc}
.param A_DWC_P  = {NP_SPLIT ? a_dwc_p  : a_dwc}
.param A_TOXE_P = {NP_SPLIT ? a_toxe_p : a_toxe}
.param A_VTH_P  = {NP_SPLIT ? a_vth_p  : a_vth}
.param A_U0_P   = {NP_SPLIT ? a_u0_p   : a_u0}
.param A_NF_P   = {NP_SPLIT ? a_nf_p   : a_nf}
.param A_VOFF_P = {NP_SPLIT ? a_voff_p : a_voff}
.param A_RDSW_P = {NP_SPLIT ? a_rdsw_p : a_rdsw}

* NFET family gains (k_<dev>_<family>_<x>)
.param k_nfet_a0_diff_cd = 0
.param k_nfet_a0_diff_damage = 0
.param k_nfet_a0_diff_eot = 0
.param k_nfet_a0_diff_act = 0
.param k_nfet_a0_diff_rc = 0
.param k_nfet_ags_diff_cd = 0
.param k_nfet_ags_diff_damage = 0
.param k_nfet_ags_diff_eot = 0
.param k_nfet_ags_diff_act = 0
.param k_nfet_ags_diff_rc = 0
.param k_nfet_b0_diff_cd = 0
.param k_nfet_b0_diff_damage = 0
.param k_nfet_b0_diff_eot = 0
.param k_nfet_b0_diff_act = 0
.param k_nfet_b0_diff_rc = 0
.param k_nfet_b1_diff_cd = 0
.param k_nfet_b1_diff_damage = 0
.param k_nfet_b1_diff_eot = 0
.param k_nfet_b1_diff_act = 0
.param k_nfet_b1_diff_rc = 0
.param k_nfet_dlc_diff_cd = {A_DLC_N}
.param k_nfet_dlc_diff_damage = 0
.param k_nfet_dlc_diff_eot = 0
.param k_nfet_dlc_diff_act = 0
.param k_nfet_dlc_diff_rc = 0
.param k_nfet_dwc_diff_cd = {A_DWC_N}
.param k_nfet_dwc_diff_damage = 0
.param k_nfet_dwc_diff_eot = 0
.param k_nfet_dwc_diff_act = 0
.param k_nfet_dwc_diff_rc = 0
.param k_nfet_eta0_diff_cd = 0
.param k_nfet_eta0_diff_damage = 0
.param k_nfet_eta0_diff_eot = 0
.param k_nfet_eta0_diff_act = 0
.param k_nfet_eta0_diff_rc = 0
.param k_nfet_k2_diff_cd = 0
.param k_nfet_k2_diff_damage = 0
.param k_nfet_k2_diff_eot = 0
.param k_nfet_k2_diff_act = 0
.param k_nfet_k2_diff_rc = 0
.param k_nfet_keta_diff_cd = 0
.param k_nfet_keta_diff_damage = 0
.param k_nfet_keta_diff_eot = 0
.param k_nfet_keta_diff_act = 0
.param k_nfet_keta_diff_rc = 0
.param k_nfet_kt1_diff_cd = 0
.param k_nfet_kt1_diff_damage = 0
.param k_nfet_kt1_diff_eot = 0
.param k_nfet_kt1_diff_act = 0
.param k_nfet_kt1_diff_rc = 0
.param k_nfet_lint_diff_cd = 0
.param k_nfet_lint_diff_damage = 0
.param k_nfet_lint_diff_eot = 0
.param k_nfet_lint_diff_act = 0
.param k_nfet_lint_diff_rc = 0
.param k_nfet_nfactor_diff_cd = 0
.param k_nfet_nfactor_diff_damage = {A_NF_N}
.param k_nfet_nfactor_diff_eot = 0
.param k_nfet_nfactor_diff_act = 0
.param k_nfet_nfactor_diff_rc = 0
.param k_nfet_overlap_mult_cd = 0
.param k_nfet_overlap_mult_damage = 0
.param k_nfet_overlap_mult_eot = 0
.param k_nfet_overlap_mult_act = 0
.param k_nfet_overlap_mult_rc = 0
.param k_nfet_pclm_diff_cd = 0
.param k_nfet_pclm_diff_damage = 0
.param k_nfet_pclm_diff_eot = 0
.param k_nfet_pclm_diff_act = 0
.param k_nfet_pclm_diff_rc = 0
.param k_nfet_pdits_diff_cd = 0
.param k_nfet_pdits_diff_damage = 0
.param k_nfet_pdits_diff_eot = 0
.param k_nfet_pdits_diff_act = 0
.param k_nfet_pdits_diff_rc = 0
.param k_nfet_pditsd_diff_cd = 0
.param k_nfet_pditsd_diff_damage = 0
.param k_nfet_pditsd_diff_eot = 0
.param k_nfet_pditsd_diff_act = 0
.param k_nfet_pditsd_diff_rc = 0
.param k_nfet_rdsw_diff_cd = 0
.param k_nfet_rdsw_diff_damage = 0
.param k_nfet_rdsw_diff_eot = 0
.param k_nfet_rdsw_diff_act = 0
.param k_nfet_rdsw_diff_rc = {A_RDSW_N}
.param k_nfet_rshn_mult_cd = 0
.param k_nfet_rshn_mult_damage = 0
.param k_nfet_rshn_mult_eot = 0
.param k_nfet_rshn_mult_act = 0
.param k_nfet_rshn_mult_rc = 0
.param k_nfet_toxe_mult_cd = 0
.param k_nfet_toxe_mult_damage = 0
.param k_nfet_toxe_mult_eot = {A_TOXE_N}
.param k_nfet_toxe_mult_act = 0
.param k_nfet_toxe_mult_rc = 0
.param k_nfet_tvoff_diff_cd = 0
.param k_nfet_tvoff_diff_damage = 0
.param k_nfet_tvoff_diff_eot = 0
.param k_nfet_tvoff_diff_act = 0
.param k_nfet_tvoff_diff_rc = 0
.param k_nfet_u0_diff_cd = 0
.param k_nfet_u0_diff_damage = {A_U0_N}
.param k_nfet_u0_diff_eot = 0
.param k_nfet_u0_diff_act = 0
.param k_nfet_u0_diff_rc = 0
.param k_nfet_ua_diff_cd = 0
.param k_nfet_ua_diff_damage = 0
.param k_nfet_ua_diff_eot = 0
.param k_nfet_ua_diff_act = 0
.param k_nfet_ua_diff_rc = 0
.param k_nfet_ub_diff_cd = 0
.param k_nfet_ub_diff_damage = 0
.param k_nfet_ub_diff_eot = 0
.param k_nfet_ub_diff_act = 0
.param k_nfet_ub_diff_rc = 0
.param k_nfet_voff_diff_cd = 0
.param k_nfet_voff_diff_damage = {A_VOFF_N}
.param k_nfet_voff_diff_eot = 0
.param k_nfet_voff_diff_act = 0
.param k_nfet_voff_diff_rc = 0
.param k_nfet_vsat_diff_cd = 0
.param k_nfet_vsat_diff_damage = 0
.param k_nfet_vsat_diff_eot = 0
.param k_nfet_vsat_diff_act = 0
.param k_nfet_vsat_diff_rc = 0
.param k_nfet_vth0_diff_cd = 0
.param k_nfet_vth0_diff_damage = 0
.param k_nfet_vth0_diff_eot = 0
.param k_nfet_vth0_diff_act = {A_VTH_N}
.param k_nfet_vth0_diff_rc = 0
.param k_nfet_wint_diff_cd = 0
.param k_nfet_wint_diff_damage = 0
.param k_nfet_wint_diff_eot = 0
.param k_nfet_wint_diff_act = 0
.param k_nfet_wint_diff_rc = 0

* PFET family gains (k_<dev>_<family>_<x>)
.param k_pfet_a0_diff_cd = 0
.param k_pfet_a0_diff_damage = 0
.param k_pfet_a0_diff_eot = 0
.param k_pfet_a0_diff_act = 0
.param k_pfet_a0_diff_rc = 0
.param k_pfet_agidl_diff_cd = 0
.param k_pfet_agidl_diff_damage = 0
.param k_pfet_agidl_diff_eot = 0
.param k_pfet_agidl_diff_act = 0
.param k_pfet_agidl_diff_rc = 0
.param k_pfet_ags_diff_cd = 0
.param k_pfet_ags_diff_damage = 0
.param k_pfet_ags_diff_eot = 0
.param k_pfet_ags_diff_act = 0
.param k_pfet_ags_diff_rc = 0
.param k_pfet_ajunction_mult_cd = 0
.param k_pfet_ajunction_mult_damage = 0
.param k_pfet_ajunction_mult_eot = 0
.param k_pfet_ajunction_mult_act = 0
.param k_pfet_ajunction_mult_rc = 0
.param k_pfet_b0_diff_cd = 0
.param k_pfet_b0_diff_damage = 0
.param k_pfet_b0_diff_eot = 0
.param k_pfet_b0_diff_act = 0
.param k_pfet_b0_diff_rc = 0
.param k_pfet_b1_diff_cd = 0
.param k_pfet_b1_diff_damage = 0
.param k_pfet_b1_diff_eot = 0
.param k_pfet_b1_diff_act = 0
.param k_pfet_b1_diff_rc = 0
.param k_pfet_bgidl_diff_cd = 0
.param k_pfet_bgidl_diff_damage = 0
.param k_pfet_bgidl_diff_eot = 0
.param k_pfet_bgidl_diff_act = 0
.param k_pfet_bgidl_diff_rc = 0
.param k_pfet_cgidl_diff_cd = 0
.param k_pfet_cgidl_diff_damage = 0
.param k_pfet_cgidl_diff_eot = 0
.param k_pfet_cgidl_diff_act = 0
.param k_pfet_cgidl_diff_rc = 0
.param k_pfet_dlc_diff_cd = {A_DLC_P}
.param k_pfet_dlc_diff_damage = 0
.param k_pfet_dlc_diff_eot = 0
.param k_pfet_dlc_diff_act = 0
.param k_pfet_dlc_diff_rc = 0
.param k_pfet_dwc_diff_cd = {A_DWC_P}
.param k_pfet_dwc_diff_damage = 0
.param k_pfet_dwc_diff_eot = 0
.param k_pfet_dwc_diff_act = 0
.param k_pfet_dwc_diff_rc = 0
.param k_pfet_eta0_diff_cd = 0
.param k_pfet_eta0_diff_damage = 0
.param k_pfet_eta0_diff_eot = 0
.param k_pfet_eta0_diff_act = 0
.param k_pfet_eta0_diff_rc = 0
.param k_pfet_k2_diff_cd = 0
.param k_pfet_k2_diff_damage = 0
.param k_pfet_k2_diff_eot = 0
.param k_pfet_k2_diff_act = 0
.param k_pfet_k2_diff_rc = 0
.param k_pfet_keta_diff_cd = 0
.param k_pfet_keta_diff_damage = 0
.param k_pfet_keta_diff_eot = 0
.param k_pfet_keta_diff_act = 0
.param k_pfet_keta_diff_rc = 0
.param k_pfet_kt1_diff_cd = 0
.param k_pfet_kt1_diff_damage = 0
.param k_pfet_kt1_diff_eot = 0
.param k_pfet_kt1_diff_act = 0
.param k_pfet_kt1_diff_rc = 0
.param k_pfet_lint_diff_cd = 0
.param k_pfet_lint_diff_damage = 0
.param k_pfet_lint_diff_eot = 0
.param k_pfet_lint_diff_act = 0
.param k_pfet_lint_diff_rc = 0
.param k_pfet_nfactor_diff_cd = 0
.param k_pfet_nfactor_diff_damage = {A_NF_P}
.param k_pfet_nfactor_diff_eot = 0
.param k_pfet_nfactor_diff_act = 0
.param k_pfet_nfactor_diff_rc = 0
.param k_pfet_overlap_mult_cd = 0
.param k_pfet_overlap_mult_damage = 0
.param k_pfet_overlap_mult_eot = 0
.param k_pfet_overlap_mult_act = 0
.param k_pfet_overlap_mult_rc = 0
.param k_pfet_pclm_diff_cd = 0
.param k_pfet_pclm_diff_damage = 0
.param k_pfet_pclm_diff_eot = 0
.param k_pfet_pclm_diff_act = 0
.param k_pfet_pclm_diff_rc = 0
.param k_pfet_pdits_diff_cd = 0
.param k_pfet_pdits_diff_damage = 0
.param k_pfet_pdits_diff_eot = 0
.param k_pfet_pdits_diff_act = 0
.param k_pfet_pdits_diff_rc = 0
.param k_pfet_pditsd_diff_cd = 0
.param k_pfet_pditsd_diff_damage = 0
.param k_pfet_pditsd_diff_eot = 0
.param k_pfet_pditsd_diff_act = 0
.param k_pfet_pditsd_diff_rc = 0
.param k_pfet_pjunction_mult_cd = 0
.param k_pfet_pjunction_mult_damage = 0
.param k_pfet_pjunction_mult_eot = 0
.param k_pfet_pjunction_mult_act = 0
.param k_pfet_pjunction_mult_rc = 0
.param k_pfet_rdsw_diff_cd = 0
.param k_pfet_rdsw_diff_damage = 0
.param k_pfet_rdsw_diff_eot = 0
.param k_pfet_rdsw_diff_act = 0
.param k_pfet_rdsw_diff_rc = {A_RDSW_P}
.param k_pfet_rshp_mult_cd = 0
.param k_pfet_rshp_mult_damage = 0
.param k_pfet_rshp_mult_eot = 0
.param k_pfet_rshp_mult_act = 0
.param k_pfet_rshp_mult_rc = 0
.param k_pfet_toxe_mult_cd = 0
.param k_pfet_toxe_mult_damage = 0
.param k_pfet_toxe_mult_eot = {A_TOXE_P}
.param k_pfet_toxe_mult_act = 0
.param k_pfet_toxe_mult_rc = 0
.param k_pfet_tvoff_diff_cd = 0
.param k_pfet_tvoff_diff_damage = 0
.param k_pfet_tvoff_diff_eot = 0
.param k_pfet_tvoff_diff_act = 0
.param k_pfet_tvoff_diff_rc = 0
.param k_pfet_u0_diff_cd = 0
.param k_pfet_u0_diff_damage = {A_U0_P}
.param k_pfet_u0_diff_eot = 0
.param k_pfet_u0_diff_act = 0
.param k_pfet_u0_diff_rc = 0
.param k_pfet_ua_diff_cd = 0
.param k_pfet_ua_diff_damage = 0
.param k_pfet_ua_diff_eot = 0
.param k_pfet_ua_diff_act = 0
.param k_pfet_ua_diff_rc = 0
.param k_pfet_ub_diff_cd = 0
.param k_pfet_ub_diff_damage = 0
.param k_pfet_ub_diff_eot = 0
.param k_pfet_ub_diff_act = 0
.param k_pfet_ub_diff_rc = 0
.param k_pfet_voff_diff_cd = 0
.param k_pfet_voff_diff_damage = {A_VOFF_P}
.param k_pfet_voff_diff_eot = 0
.param k_pfet_voff_diff_act = 0
.param k_pfet_voff_diff_rc = 0
.param k_pfet_vsat_diff_cd = 0
.param k_pfet_vsat_diff_damage = 0
.param k_pfet_vsat_diff_eot = 0
.param k_pfet_vsat_diff_act = 0
.param k_pfet_vsat_diff_rc = 0
.param k_pfet_vth0_diff_cd = 0
.param k_pfet_vth0_diff_damage = 0
.param k_pfet_vth0_diff_eot = 0
.param k_pfet_vth0_diff_act = {A_VTH_P}
.param k_pfet_vth0_diff_rc = 0
.param k_pfet_wint_diff_cd = 0
.param k_pfet_wint_diff_damage = 0
.param k_pfet_wint_diff_eot = 0
.param k_pfet_wint_diff_act = 0
.param k_pfet_wint_diff_rc = 0

* Full wafer variable mapping equations
* NFET equations
.param sky130_fd_pr__nfet_01v8__dlc_diff = {sky130_fd_pr__nfet_01v8__dlc_diff + k_nfet_dlc_diff_cd*X_cd + k_nfet_dlc_diff_damage*X_damage + k_nfet_dlc_diff_eot*X_eot + k_nfet_dlc_diff_act*X_act + k_nfet_dlc_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__dwc_diff = {sky130_fd_pr__nfet_01v8__dwc_diff + k_nfet_dwc_diff_cd*X_cd + k_nfet_dwc_diff_damage*X_damage + k_nfet_dwc_diff_eot*X_eot + k_nfet_dwc_diff_act*X_act + k_nfet_dwc_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__lint_diff = {sky130_fd_pr__nfet_01v8__lint_diff + k_nfet_lint_diff_cd*X_cd + k_nfet_lint_diff_damage*X_damage + k_nfet_lint_diff_eot*X_eot + k_nfet_lint_diff_act*X_act + k_nfet_lint_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__overlap_mult = {sky130_fd_pr__nfet_01v8__overlap_mult*(1 + k_nfet_overlap_mult_cd*X_cd + k_nfet_overlap_mult_damage*X_damage + k_nfet_overlap_mult_eot*X_eot + k_nfet_overlap_mult_act*X_act + k_nfet_overlap_mult_rc*X_rc)}
.param sky130_fd_pr__nfet_01v8__rshn_mult = {sky130_fd_pr__nfet_01v8__rshn_mult*(1 + k_nfet_rshn_mult_cd*X_cd + k_nfet_rshn_mult_damage*X_damage + k_nfet_rshn_mult_eot*X_eot + k_nfet_rshn_mult_act*X_act + k_nfet_rshn_mult_rc*X_rc)}
.param sky130_fd_pr__nfet_01v8__toxe_mult = {sky130_fd_pr__nfet_01v8__toxe_mult*(1 + k_nfet_toxe_mult_cd*X_cd + k_nfet_toxe_mult_damage*X_damage + k_nfet_toxe_mult_eot*X_eot + k_nfet_toxe_mult_act*X_act + k_nfet_toxe_mult_rc*X_rc)}
.param sky130_fd_pr__nfet_01v8__wint_diff = {sky130_fd_pr__nfet_01v8__wint_diff + k_nfet_wint_diff_cd*X_cd + k_nfet_wint_diff_damage*X_damage + k_nfet_wint_diff_eot*X_eot + k_nfet_wint_diff_act*X_act + k_nfet_wint_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_0 = {sky130_fd_pr__nfet_01v8__a0_diff_0 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_1 = {sky130_fd_pr__nfet_01v8__a0_diff_1 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_10 = {sky130_fd_pr__nfet_01v8__a0_diff_10 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_11 = {sky130_fd_pr__nfet_01v8__a0_diff_11 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_12 = {sky130_fd_pr__nfet_01v8__a0_diff_12 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_13 = {sky130_fd_pr__nfet_01v8__a0_diff_13 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_14 = {sky130_fd_pr__nfet_01v8__a0_diff_14 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_15 = {sky130_fd_pr__nfet_01v8__a0_diff_15 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_16 = {sky130_fd_pr__nfet_01v8__a0_diff_16 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_17 = {sky130_fd_pr__nfet_01v8__a0_diff_17 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_18 = {sky130_fd_pr__nfet_01v8__a0_diff_18 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_19 = {sky130_fd_pr__nfet_01v8__a0_diff_19 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_2 = {sky130_fd_pr__nfet_01v8__a0_diff_2 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_20 = {sky130_fd_pr__nfet_01v8__a0_diff_20 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_21 = {sky130_fd_pr__nfet_01v8__a0_diff_21 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_22 = {sky130_fd_pr__nfet_01v8__a0_diff_22 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_23 = {sky130_fd_pr__nfet_01v8__a0_diff_23 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_24 = {sky130_fd_pr__nfet_01v8__a0_diff_24 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_25 = {sky130_fd_pr__nfet_01v8__a0_diff_25 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_26 = {sky130_fd_pr__nfet_01v8__a0_diff_26 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_27 = {sky130_fd_pr__nfet_01v8__a0_diff_27 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_28 = {sky130_fd_pr__nfet_01v8__a0_diff_28 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_29 = {sky130_fd_pr__nfet_01v8__a0_diff_29 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_3 = {sky130_fd_pr__nfet_01v8__a0_diff_3 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_30 = {sky130_fd_pr__nfet_01v8__a0_diff_30 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_31 = {sky130_fd_pr__nfet_01v8__a0_diff_31 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_32 = {sky130_fd_pr__nfet_01v8__a0_diff_32 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_33 = {sky130_fd_pr__nfet_01v8__a0_diff_33 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_34 = {sky130_fd_pr__nfet_01v8__a0_diff_34 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_35 = {sky130_fd_pr__nfet_01v8__a0_diff_35 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_36 = {sky130_fd_pr__nfet_01v8__a0_diff_36 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_37 = {sky130_fd_pr__nfet_01v8__a0_diff_37 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_38 = {sky130_fd_pr__nfet_01v8__a0_diff_38 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_39 = {sky130_fd_pr__nfet_01v8__a0_diff_39 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_4 = {sky130_fd_pr__nfet_01v8__a0_diff_4 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_40 = {sky130_fd_pr__nfet_01v8__a0_diff_40 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_41 = {sky130_fd_pr__nfet_01v8__a0_diff_41 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_42 = {sky130_fd_pr__nfet_01v8__a0_diff_42 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_43 = {sky130_fd_pr__nfet_01v8__a0_diff_43 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_44 = {sky130_fd_pr__nfet_01v8__a0_diff_44 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_45 = {sky130_fd_pr__nfet_01v8__a0_diff_45 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_46 = {sky130_fd_pr__nfet_01v8__a0_diff_46 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_47 = {sky130_fd_pr__nfet_01v8__a0_diff_47 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_48 = {sky130_fd_pr__nfet_01v8__a0_diff_48 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_49 = {sky130_fd_pr__nfet_01v8__a0_diff_49 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_5 = {sky130_fd_pr__nfet_01v8__a0_diff_5 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_50 = {sky130_fd_pr__nfet_01v8__a0_diff_50 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_51 = {sky130_fd_pr__nfet_01v8__a0_diff_51 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_52 = {sky130_fd_pr__nfet_01v8__a0_diff_52 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_53 = {sky130_fd_pr__nfet_01v8__a0_diff_53 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_54 = {sky130_fd_pr__nfet_01v8__a0_diff_54 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_55 = {sky130_fd_pr__nfet_01v8__a0_diff_55 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_56 = {sky130_fd_pr__nfet_01v8__a0_diff_56 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_57 = {sky130_fd_pr__nfet_01v8__a0_diff_57 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_58 = {sky130_fd_pr__nfet_01v8__a0_diff_58 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_59 = {sky130_fd_pr__nfet_01v8__a0_diff_59 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_6 = {sky130_fd_pr__nfet_01v8__a0_diff_6 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_60 = {sky130_fd_pr__nfet_01v8__a0_diff_60 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_61 = {sky130_fd_pr__nfet_01v8__a0_diff_61 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_62 = {sky130_fd_pr__nfet_01v8__a0_diff_62 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_7 = {sky130_fd_pr__nfet_01v8__a0_diff_7 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_8 = {sky130_fd_pr__nfet_01v8__a0_diff_8 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__a0_diff_9 = {sky130_fd_pr__nfet_01v8__a0_diff_9 + k_nfet_a0_diff_cd*X_cd + k_nfet_a0_diff_damage*X_damage + k_nfet_a0_diff_eot*X_eot + k_nfet_a0_diff_act*X_act + k_nfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_0 = {sky130_fd_pr__nfet_01v8__ags_diff_0 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_1 = {sky130_fd_pr__nfet_01v8__ags_diff_1 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_10 = {sky130_fd_pr__nfet_01v8__ags_diff_10 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_11 = {sky130_fd_pr__nfet_01v8__ags_diff_11 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_12 = {sky130_fd_pr__nfet_01v8__ags_diff_12 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_13 = {sky130_fd_pr__nfet_01v8__ags_diff_13 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_14 = {sky130_fd_pr__nfet_01v8__ags_diff_14 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_15 = {sky130_fd_pr__nfet_01v8__ags_diff_15 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_16 = {sky130_fd_pr__nfet_01v8__ags_diff_16 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_17 = {sky130_fd_pr__nfet_01v8__ags_diff_17 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_18 = {sky130_fd_pr__nfet_01v8__ags_diff_18 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_19 = {sky130_fd_pr__nfet_01v8__ags_diff_19 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_2 = {sky130_fd_pr__nfet_01v8__ags_diff_2 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_20 = {sky130_fd_pr__nfet_01v8__ags_diff_20 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_21 = {sky130_fd_pr__nfet_01v8__ags_diff_21 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_22 = {sky130_fd_pr__nfet_01v8__ags_diff_22 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_23 = {sky130_fd_pr__nfet_01v8__ags_diff_23 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_24 = {sky130_fd_pr__nfet_01v8__ags_diff_24 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_25 = {sky130_fd_pr__nfet_01v8__ags_diff_25 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_26 = {sky130_fd_pr__nfet_01v8__ags_diff_26 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_27 = {sky130_fd_pr__nfet_01v8__ags_diff_27 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_28 = {sky130_fd_pr__nfet_01v8__ags_diff_28 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_29 = {sky130_fd_pr__nfet_01v8__ags_diff_29 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_3 = {sky130_fd_pr__nfet_01v8__ags_diff_3 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_30 = {sky130_fd_pr__nfet_01v8__ags_diff_30 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_31 = {sky130_fd_pr__nfet_01v8__ags_diff_31 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_32 = {sky130_fd_pr__nfet_01v8__ags_diff_32 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_33 = {sky130_fd_pr__nfet_01v8__ags_diff_33 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_34 = {sky130_fd_pr__nfet_01v8__ags_diff_34 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_35 = {sky130_fd_pr__nfet_01v8__ags_diff_35 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_36 = {sky130_fd_pr__nfet_01v8__ags_diff_36 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_37 = {sky130_fd_pr__nfet_01v8__ags_diff_37 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_38 = {sky130_fd_pr__nfet_01v8__ags_diff_38 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_39 = {sky130_fd_pr__nfet_01v8__ags_diff_39 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_4 = {sky130_fd_pr__nfet_01v8__ags_diff_4 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_40 = {sky130_fd_pr__nfet_01v8__ags_diff_40 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_41 = {sky130_fd_pr__nfet_01v8__ags_diff_41 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_42 = {sky130_fd_pr__nfet_01v8__ags_diff_42 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_43 = {sky130_fd_pr__nfet_01v8__ags_diff_43 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_44 = {sky130_fd_pr__nfet_01v8__ags_diff_44 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_45 = {sky130_fd_pr__nfet_01v8__ags_diff_45 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_46 = {sky130_fd_pr__nfet_01v8__ags_diff_46 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_47 = {sky130_fd_pr__nfet_01v8__ags_diff_47 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_48 = {sky130_fd_pr__nfet_01v8__ags_diff_48 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_49 = {sky130_fd_pr__nfet_01v8__ags_diff_49 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_5 = {sky130_fd_pr__nfet_01v8__ags_diff_5 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_50 = {sky130_fd_pr__nfet_01v8__ags_diff_50 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_51 = {sky130_fd_pr__nfet_01v8__ags_diff_51 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_52 = {sky130_fd_pr__nfet_01v8__ags_diff_52 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_53 = {sky130_fd_pr__nfet_01v8__ags_diff_53 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_54 = {sky130_fd_pr__nfet_01v8__ags_diff_54 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_55 = {sky130_fd_pr__nfet_01v8__ags_diff_55 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_56 = {sky130_fd_pr__nfet_01v8__ags_diff_56 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_57 = {sky130_fd_pr__nfet_01v8__ags_diff_57 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_58 = {sky130_fd_pr__nfet_01v8__ags_diff_58 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_59 = {sky130_fd_pr__nfet_01v8__ags_diff_59 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_6 = {sky130_fd_pr__nfet_01v8__ags_diff_6 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_60 = {sky130_fd_pr__nfet_01v8__ags_diff_60 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_61 = {sky130_fd_pr__nfet_01v8__ags_diff_61 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_62 = {sky130_fd_pr__nfet_01v8__ags_diff_62 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_7 = {sky130_fd_pr__nfet_01v8__ags_diff_7 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_8 = {sky130_fd_pr__nfet_01v8__ags_diff_8 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ags_diff_9 = {sky130_fd_pr__nfet_01v8__ags_diff_9 + k_nfet_ags_diff_cd*X_cd + k_nfet_ags_diff_damage*X_damage + k_nfet_ags_diff_eot*X_eot + k_nfet_ags_diff_act*X_act + k_nfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_0 = {sky130_fd_pr__nfet_01v8__b0_diff_0 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_1 = {sky130_fd_pr__nfet_01v8__b0_diff_1 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_10 = {sky130_fd_pr__nfet_01v8__b0_diff_10 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_11 = {sky130_fd_pr__nfet_01v8__b0_diff_11 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_12 = {sky130_fd_pr__nfet_01v8__b0_diff_12 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_13 = {sky130_fd_pr__nfet_01v8__b0_diff_13 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_14 = {sky130_fd_pr__nfet_01v8__b0_diff_14 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_15 = {sky130_fd_pr__nfet_01v8__b0_diff_15 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_16 = {sky130_fd_pr__nfet_01v8__b0_diff_16 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_17 = {sky130_fd_pr__nfet_01v8__b0_diff_17 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_18 = {sky130_fd_pr__nfet_01v8__b0_diff_18 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_19 = {sky130_fd_pr__nfet_01v8__b0_diff_19 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_2 = {sky130_fd_pr__nfet_01v8__b0_diff_2 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_20 = {sky130_fd_pr__nfet_01v8__b0_diff_20 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_21 = {sky130_fd_pr__nfet_01v8__b0_diff_21 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_22 = {sky130_fd_pr__nfet_01v8__b0_diff_22 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_23 = {sky130_fd_pr__nfet_01v8__b0_diff_23 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_24 = {sky130_fd_pr__nfet_01v8__b0_diff_24 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_25 = {sky130_fd_pr__nfet_01v8__b0_diff_25 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_26 = {sky130_fd_pr__nfet_01v8__b0_diff_26 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_27 = {sky130_fd_pr__nfet_01v8__b0_diff_27 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_28 = {sky130_fd_pr__nfet_01v8__b0_diff_28 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_29 = {sky130_fd_pr__nfet_01v8__b0_diff_29 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_3 = {sky130_fd_pr__nfet_01v8__b0_diff_3 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_30 = {sky130_fd_pr__nfet_01v8__b0_diff_30 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_31 = {sky130_fd_pr__nfet_01v8__b0_diff_31 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_32 = {sky130_fd_pr__nfet_01v8__b0_diff_32 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_33 = {sky130_fd_pr__nfet_01v8__b0_diff_33 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_34 = {sky130_fd_pr__nfet_01v8__b0_diff_34 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_35 = {sky130_fd_pr__nfet_01v8__b0_diff_35 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_36 = {sky130_fd_pr__nfet_01v8__b0_diff_36 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_37 = {sky130_fd_pr__nfet_01v8__b0_diff_37 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_38 = {sky130_fd_pr__nfet_01v8__b0_diff_38 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_39 = {sky130_fd_pr__nfet_01v8__b0_diff_39 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_4 = {sky130_fd_pr__nfet_01v8__b0_diff_4 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_40 = {sky130_fd_pr__nfet_01v8__b0_diff_40 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_41 = {sky130_fd_pr__nfet_01v8__b0_diff_41 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_42 = {sky130_fd_pr__nfet_01v8__b0_diff_42 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_43 = {sky130_fd_pr__nfet_01v8__b0_diff_43 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_44 = {sky130_fd_pr__nfet_01v8__b0_diff_44 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_45 = {sky130_fd_pr__nfet_01v8__b0_diff_45 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_46 = {sky130_fd_pr__nfet_01v8__b0_diff_46 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_47 = {sky130_fd_pr__nfet_01v8__b0_diff_47 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_48 = {sky130_fd_pr__nfet_01v8__b0_diff_48 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_49 = {sky130_fd_pr__nfet_01v8__b0_diff_49 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_5 = {sky130_fd_pr__nfet_01v8__b0_diff_5 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_50 = {sky130_fd_pr__nfet_01v8__b0_diff_50 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_51 = {sky130_fd_pr__nfet_01v8__b0_diff_51 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_52 = {sky130_fd_pr__nfet_01v8__b0_diff_52 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_53 = {sky130_fd_pr__nfet_01v8__b0_diff_53 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_54 = {sky130_fd_pr__nfet_01v8__b0_diff_54 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_55 = {sky130_fd_pr__nfet_01v8__b0_diff_55 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_56 = {sky130_fd_pr__nfet_01v8__b0_diff_56 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_57 = {sky130_fd_pr__nfet_01v8__b0_diff_57 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_58 = {sky130_fd_pr__nfet_01v8__b0_diff_58 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_59 = {sky130_fd_pr__nfet_01v8__b0_diff_59 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_6 = {sky130_fd_pr__nfet_01v8__b0_diff_6 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_60 = {sky130_fd_pr__nfet_01v8__b0_diff_60 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_61 = {sky130_fd_pr__nfet_01v8__b0_diff_61 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_62 = {sky130_fd_pr__nfet_01v8__b0_diff_62 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_7 = {sky130_fd_pr__nfet_01v8__b0_diff_7 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_8 = {sky130_fd_pr__nfet_01v8__b0_diff_8 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b0_diff_9 = {sky130_fd_pr__nfet_01v8__b0_diff_9 + k_nfet_b0_diff_cd*X_cd + k_nfet_b0_diff_damage*X_damage + k_nfet_b0_diff_eot*X_eot + k_nfet_b0_diff_act*X_act + k_nfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_0 = {sky130_fd_pr__nfet_01v8__b1_diff_0 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_1 = {sky130_fd_pr__nfet_01v8__b1_diff_1 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_10 = {sky130_fd_pr__nfet_01v8__b1_diff_10 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_11 = {sky130_fd_pr__nfet_01v8__b1_diff_11 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_12 = {sky130_fd_pr__nfet_01v8__b1_diff_12 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_13 = {sky130_fd_pr__nfet_01v8__b1_diff_13 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_14 = {sky130_fd_pr__nfet_01v8__b1_diff_14 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_15 = {sky130_fd_pr__nfet_01v8__b1_diff_15 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_16 = {sky130_fd_pr__nfet_01v8__b1_diff_16 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_17 = {sky130_fd_pr__nfet_01v8__b1_diff_17 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_18 = {sky130_fd_pr__nfet_01v8__b1_diff_18 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_19 = {sky130_fd_pr__nfet_01v8__b1_diff_19 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_2 = {sky130_fd_pr__nfet_01v8__b1_diff_2 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_20 = {sky130_fd_pr__nfet_01v8__b1_diff_20 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_21 = {sky130_fd_pr__nfet_01v8__b1_diff_21 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_22 = {sky130_fd_pr__nfet_01v8__b1_diff_22 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_23 = {sky130_fd_pr__nfet_01v8__b1_diff_23 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_24 = {sky130_fd_pr__nfet_01v8__b1_diff_24 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_25 = {sky130_fd_pr__nfet_01v8__b1_diff_25 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_26 = {sky130_fd_pr__nfet_01v8__b1_diff_26 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_27 = {sky130_fd_pr__nfet_01v8__b1_diff_27 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_28 = {sky130_fd_pr__nfet_01v8__b1_diff_28 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_29 = {sky130_fd_pr__nfet_01v8__b1_diff_29 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_3 = {sky130_fd_pr__nfet_01v8__b1_diff_3 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_30 = {sky130_fd_pr__nfet_01v8__b1_diff_30 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_31 = {sky130_fd_pr__nfet_01v8__b1_diff_31 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_32 = {sky130_fd_pr__nfet_01v8__b1_diff_32 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_33 = {sky130_fd_pr__nfet_01v8__b1_diff_33 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_34 = {sky130_fd_pr__nfet_01v8__b1_diff_34 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_35 = {sky130_fd_pr__nfet_01v8__b1_diff_35 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_36 = {sky130_fd_pr__nfet_01v8__b1_diff_36 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_37 = {sky130_fd_pr__nfet_01v8__b1_diff_37 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_38 = {sky130_fd_pr__nfet_01v8__b1_diff_38 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_39 = {sky130_fd_pr__nfet_01v8__b1_diff_39 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_4 = {sky130_fd_pr__nfet_01v8__b1_diff_4 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_40 = {sky130_fd_pr__nfet_01v8__b1_diff_40 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_41 = {sky130_fd_pr__nfet_01v8__b1_diff_41 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_42 = {sky130_fd_pr__nfet_01v8__b1_diff_42 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_43 = {sky130_fd_pr__nfet_01v8__b1_diff_43 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_44 = {sky130_fd_pr__nfet_01v8__b1_diff_44 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_45 = {sky130_fd_pr__nfet_01v8__b1_diff_45 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_46 = {sky130_fd_pr__nfet_01v8__b1_diff_46 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_47 = {sky130_fd_pr__nfet_01v8__b1_diff_47 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_48 = {sky130_fd_pr__nfet_01v8__b1_diff_48 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_49 = {sky130_fd_pr__nfet_01v8__b1_diff_49 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_5 = {sky130_fd_pr__nfet_01v8__b1_diff_5 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_50 = {sky130_fd_pr__nfet_01v8__b1_diff_50 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_51 = {sky130_fd_pr__nfet_01v8__b1_diff_51 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_52 = {sky130_fd_pr__nfet_01v8__b1_diff_52 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_53 = {sky130_fd_pr__nfet_01v8__b1_diff_53 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_54 = {sky130_fd_pr__nfet_01v8__b1_diff_54 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_55 = {sky130_fd_pr__nfet_01v8__b1_diff_55 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_56 = {sky130_fd_pr__nfet_01v8__b1_diff_56 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_57 = {sky130_fd_pr__nfet_01v8__b1_diff_57 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_58 = {sky130_fd_pr__nfet_01v8__b1_diff_58 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_59 = {sky130_fd_pr__nfet_01v8__b1_diff_59 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_6 = {sky130_fd_pr__nfet_01v8__b1_diff_6 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_60 = {sky130_fd_pr__nfet_01v8__b1_diff_60 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_61 = {sky130_fd_pr__nfet_01v8__b1_diff_61 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_62 = {sky130_fd_pr__nfet_01v8__b1_diff_62 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_7 = {sky130_fd_pr__nfet_01v8__b1_diff_7 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_8 = {sky130_fd_pr__nfet_01v8__b1_diff_8 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__b1_diff_9 = {sky130_fd_pr__nfet_01v8__b1_diff_9 + k_nfet_b1_diff_cd*X_cd + k_nfet_b1_diff_damage*X_damage + k_nfet_b1_diff_eot*X_eot + k_nfet_b1_diff_act*X_act + k_nfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_0 = {sky130_fd_pr__nfet_01v8__eta0_diff_0 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_1 = {sky130_fd_pr__nfet_01v8__eta0_diff_1 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_10 = {sky130_fd_pr__nfet_01v8__eta0_diff_10 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_11 = {sky130_fd_pr__nfet_01v8__eta0_diff_11 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_12 = {sky130_fd_pr__nfet_01v8__eta0_diff_12 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_13 = {sky130_fd_pr__nfet_01v8__eta0_diff_13 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_14 = {sky130_fd_pr__nfet_01v8__eta0_diff_14 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_15 = {sky130_fd_pr__nfet_01v8__eta0_diff_15 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_16 = {sky130_fd_pr__nfet_01v8__eta0_diff_16 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_17 = {sky130_fd_pr__nfet_01v8__eta0_diff_17 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_18 = {sky130_fd_pr__nfet_01v8__eta0_diff_18 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_19 = {sky130_fd_pr__nfet_01v8__eta0_diff_19 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_2 = {sky130_fd_pr__nfet_01v8__eta0_diff_2 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_20 = {sky130_fd_pr__nfet_01v8__eta0_diff_20 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_21 = {sky130_fd_pr__nfet_01v8__eta0_diff_21 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_22 = {sky130_fd_pr__nfet_01v8__eta0_diff_22 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_23 = {sky130_fd_pr__nfet_01v8__eta0_diff_23 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_24 = {sky130_fd_pr__nfet_01v8__eta0_diff_24 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_25 = {sky130_fd_pr__nfet_01v8__eta0_diff_25 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_26 = {sky130_fd_pr__nfet_01v8__eta0_diff_26 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_27 = {sky130_fd_pr__nfet_01v8__eta0_diff_27 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_28 = {sky130_fd_pr__nfet_01v8__eta0_diff_28 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_29 = {sky130_fd_pr__nfet_01v8__eta0_diff_29 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_3 = {sky130_fd_pr__nfet_01v8__eta0_diff_3 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_30 = {sky130_fd_pr__nfet_01v8__eta0_diff_30 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_31 = {sky130_fd_pr__nfet_01v8__eta0_diff_31 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_32 = {sky130_fd_pr__nfet_01v8__eta0_diff_32 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_33 = {sky130_fd_pr__nfet_01v8__eta0_diff_33 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_34 = {sky130_fd_pr__nfet_01v8__eta0_diff_34 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_35 = {sky130_fd_pr__nfet_01v8__eta0_diff_35 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_36 = {sky130_fd_pr__nfet_01v8__eta0_diff_36 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_37 = {sky130_fd_pr__nfet_01v8__eta0_diff_37 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_38 = {sky130_fd_pr__nfet_01v8__eta0_diff_38 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_39 = {sky130_fd_pr__nfet_01v8__eta0_diff_39 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_4 = {sky130_fd_pr__nfet_01v8__eta0_diff_4 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_40 = {sky130_fd_pr__nfet_01v8__eta0_diff_40 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_41 = {sky130_fd_pr__nfet_01v8__eta0_diff_41 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_42 = {sky130_fd_pr__nfet_01v8__eta0_diff_42 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_43 = {sky130_fd_pr__nfet_01v8__eta0_diff_43 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_44 = {sky130_fd_pr__nfet_01v8__eta0_diff_44 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_45 = {sky130_fd_pr__nfet_01v8__eta0_diff_45 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_46 = {sky130_fd_pr__nfet_01v8__eta0_diff_46 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_47 = {sky130_fd_pr__nfet_01v8__eta0_diff_47 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_48 = {sky130_fd_pr__nfet_01v8__eta0_diff_48 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_49 = {sky130_fd_pr__nfet_01v8__eta0_diff_49 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_5 = {sky130_fd_pr__nfet_01v8__eta0_diff_5 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_50 = {sky130_fd_pr__nfet_01v8__eta0_diff_50 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_51 = {sky130_fd_pr__nfet_01v8__eta0_diff_51 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_52 = {sky130_fd_pr__nfet_01v8__eta0_diff_52 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_53 = {sky130_fd_pr__nfet_01v8__eta0_diff_53 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_54 = {sky130_fd_pr__nfet_01v8__eta0_diff_54 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_55 = {sky130_fd_pr__nfet_01v8__eta0_diff_55 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_56 = {sky130_fd_pr__nfet_01v8__eta0_diff_56 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_57 = {sky130_fd_pr__nfet_01v8__eta0_diff_57 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_58 = {sky130_fd_pr__nfet_01v8__eta0_diff_58 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_59 = {sky130_fd_pr__nfet_01v8__eta0_diff_59 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_6 = {sky130_fd_pr__nfet_01v8__eta0_diff_6 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_60 = {sky130_fd_pr__nfet_01v8__eta0_diff_60 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_61 = {sky130_fd_pr__nfet_01v8__eta0_diff_61 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_62 = {sky130_fd_pr__nfet_01v8__eta0_diff_62 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_7 = {sky130_fd_pr__nfet_01v8__eta0_diff_7 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_8 = {sky130_fd_pr__nfet_01v8__eta0_diff_8 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__eta0_diff_9 = {sky130_fd_pr__nfet_01v8__eta0_diff_9 + k_nfet_eta0_diff_cd*X_cd + k_nfet_eta0_diff_damage*X_damage + k_nfet_eta0_diff_eot*X_eot + k_nfet_eta0_diff_act*X_act + k_nfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_0 = {sky130_fd_pr__nfet_01v8__k2_diff_0 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_1 = {sky130_fd_pr__nfet_01v8__k2_diff_1 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_10 = {sky130_fd_pr__nfet_01v8__k2_diff_10 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_11 = {sky130_fd_pr__nfet_01v8__k2_diff_11 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_12 = {sky130_fd_pr__nfet_01v8__k2_diff_12 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_13 = {sky130_fd_pr__nfet_01v8__k2_diff_13 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_14 = {sky130_fd_pr__nfet_01v8__k2_diff_14 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_15 = {sky130_fd_pr__nfet_01v8__k2_diff_15 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_16 = {sky130_fd_pr__nfet_01v8__k2_diff_16 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_17 = {sky130_fd_pr__nfet_01v8__k2_diff_17 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_18 = {sky130_fd_pr__nfet_01v8__k2_diff_18 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_19 = {sky130_fd_pr__nfet_01v8__k2_diff_19 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_2 = {sky130_fd_pr__nfet_01v8__k2_diff_2 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_20 = {sky130_fd_pr__nfet_01v8__k2_diff_20 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_21 = {sky130_fd_pr__nfet_01v8__k2_diff_21 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_22 = {sky130_fd_pr__nfet_01v8__k2_diff_22 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_23 = {sky130_fd_pr__nfet_01v8__k2_diff_23 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_24 = {sky130_fd_pr__nfet_01v8__k2_diff_24 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_25 = {sky130_fd_pr__nfet_01v8__k2_diff_25 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_26 = {sky130_fd_pr__nfet_01v8__k2_diff_26 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_27 = {sky130_fd_pr__nfet_01v8__k2_diff_27 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_28 = {sky130_fd_pr__nfet_01v8__k2_diff_28 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_29 = {sky130_fd_pr__nfet_01v8__k2_diff_29 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_3 = {sky130_fd_pr__nfet_01v8__k2_diff_3 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_30 = {sky130_fd_pr__nfet_01v8__k2_diff_30 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_31 = {sky130_fd_pr__nfet_01v8__k2_diff_31 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_32 = {sky130_fd_pr__nfet_01v8__k2_diff_32 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_33 = {sky130_fd_pr__nfet_01v8__k2_diff_33 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_34 = {sky130_fd_pr__nfet_01v8__k2_diff_34 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_35 = {sky130_fd_pr__nfet_01v8__k2_diff_35 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_36 = {sky130_fd_pr__nfet_01v8__k2_diff_36 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_37 = {sky130_fd_pr__nfet_01v8__k2_diff_37 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_38 = {sky130_fd_pr__nfet_01v8__k2_diff_38 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_39 = {sky130_fd_pr__nfet_01v8__k2_diff_39 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_4 = {sky130_fd_pr__nfet_01v8__k2_diff_4 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_40 = {sky130_fd_pr__nfet_01v8__k2_diff_40 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_41 = {sky130_fd_pr__nfet_01v8__k2_diff_41 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_42 = {sky130_fd_pr__nfet_01v8__k2_diff_42 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_43 = {sky130_fd_pr__nfet_01v8__k2_diff_43 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_44 = {sky130_fd_pr__nfet_01v8__k2_diff_44 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_45 = {sky130_fd_pr__nfet_01v8__k2_diff_45 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_46 = {sky130_fd_pr__nfet_01v8__k2_diff_46 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_47 = {sky130_fd_pr__nfet_01v8__k2_diff_47 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_48 = {sky130_fd_pr__nfet_01v8__k2_diff_48 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_49 = {sky130_fd_pr__nfet_01v8__k2_diff_49 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_5 = {sky130_fd_pr__nfet_01v8__k2_diff_5 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_50 = {sky130_fd_pr__nfet_01v8__k2_diff_50 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_51 = {sky130_fd_pr__nfet_01v8__k2_diff_51 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_52 = {sky130_fd_pr__nfet_01v8__k2_diff_52 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_53 = {sky130_fd_pr__nfet_01v8__k2_diff_53 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_54 = {sky130_fd_pr__nfet_01v8__k2_diff_54 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_55 = {sky130_fd_pr__nfet_01v8__k2_diff_55 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_56 = {sky130_fd_pr__nfet_01v8__k2_diff_56 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_57 = {sky130_fd_pr__nfet_01v8__k2_diff_57 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_58 = {sky130_fd_pr__nfet_01v8__k2_diff_58 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_59 = {sky130_fd_pr__nfet_01v8__k2_diff_59 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_6 = {sky130_fd_pr__nfet_01v8__k2_diff_6 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_60 = {sky130_fd_pr__nfet_01v8__k2_diff_60 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_61 = {sky130_fd_pr__nfet_01v8__k2_diff_61 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_62 = {sky130_fd_pr__nfet_01v8__k2_diff_62 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_7 = {sky130_fd_pr__nfet_01v8__k2_diff_7 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_8 = {sky130_fd_pr__nfet_01v8__k2_diff_8 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__k2_diff_9 = {sky130_fd_pr__nfet_01v8__k2_diff_9 + k_nfet_k2_diff_cd*X_cd + k_nfet_k2_diff_damage*X_damage + k_nfet_k2_diff_eot*X_eot + k_nfet_k2_diff_act*X_act + k_nfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_0 = {sky130_fd_pr__nfet_01v8__keta_diff_0 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_1 = {sky130_fd_pr__nfet_01v8__keta_diff_1 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_10 = {sky130_fd_pr__nfet_01v8__keta_diff_10 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_11 = {sky130_fd_pr__nfet_01v8__keta_diff_11 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_12 = {sky130_fd_pr__nfet_01v8__keta_diff_12 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_13 = {sky130_fd_pr__nfet_01v8__keta_diff_13 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_14 = {sky130_fd_pr__nfet_01v8__keta_diff_14 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_15 = {sky130_fd_pr__nfet_01v8__keta_diff_15 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_16 = {sky130_fd_pr__nfet_01v8__keta_diff_16 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_17 = {sky130_fd_pr__nfet_01v8__keta_diff_17 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_18 = {sky130_fd_pr__nfet_01v8__keta_diff_18 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_19 = {sky130_fd_pr__nfet_01v8__keta_diff_19 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_2 = {sky130_fd_pr__nfet_01v8__keta_diff_2 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_20 = {sky130_fd_pr__nfet_01v8__keta_diff_20 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_21 = {sky130_fd_pr__nfet_01v8__keta_diff_21 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_22 = {sky130_fd_pr__nfet_01v8__keta_diff_22 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_23 = {sky130_fd_pr__nfet_01v8__keta_diff_23 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_24 = {sky130_fd_pr__nfet_01v8__keta_diff_24 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_25 = {sky130_fd_pr__nfet_01v8__keta_diff_25 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_26 = {sky130_fd_pr__nfet_01v8__keta_diff_26 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_27 = {sky130_fd_pr__nfet_01v8__keta_diff_27 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_28 = {sky130_fd_pr__nfet_01v8__keta_diff_28 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_29 = {sky130_fd_pr__nfet_01v8__keta_diff_29 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_3 = {sky130_fd_pr__nfet_01v8__keta_diff_3 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_30 = {sky130_fd_pr__nfet_01v8__keta_diff_30 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_31 = {sky130_fd_pr__nfet_01v8__keta_diff_31 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_32 = {sky130_fd_pr__nfet_01v8__keta_diff_32 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_33 = {sky130_fd_pr__nfet_01v8__keta_diff_33 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_34 = {sky130_fd_pr__nfet_01v8__keta_diff_34 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_35 = {sky130_fd_pr__nfet_01v8__keta_diff_35 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_36 = {sky130_fd_pr__nfet_01v8__keta_diff_36 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_37 = {sky130_fd_pr__nfet_01v8__keta_diff_37 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_38 = {sky130_fd_pr__nfet_01v8__keta_diff_38 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_39 = {sky130_fd_pr__nfet_01v8__keta_diff_39 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_4 = {sky130_fd_pr__nfet_01v8__keta_diff_4 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_40 = {sky130_fd_pr__nfet_01v8__keta_diff_40 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_41 = {sky130_fd_pr__nfet_01v8__keta_diff_41 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_42 = {sky130_fd_pr__nfet_01v8__keta_diff_42 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_43 = {sky130_fd_pr__nfet_01v8__keta_diff_43 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_44 = {sky130_fd_pr__nfet_01v8__keta_diff_44 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_45 = {sky130_fd_pr__nfet_01v8__keta_diff_45 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_46 = {sky130_fd_pr__nfet_01v8__keta_diff_46 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_47 = {sky130_fd_pr__nfet_01v8__keta_diff_47 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_48 = {sky130_fd_pr__nfet_01v8__keta_diff_48 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_49 = {sky130_fd_pr__nfet_01v8__keta_diff_49 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_5 = {sky130_fd_pr__nfet_01v8__keta_diff_5 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_50 = {sky130_fd_pr__nfet_01v8__keta_diff_50 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_51 = {sky130_fd_pr__nfet_01v8__keta_diff_51 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_52 = {sky130_fd_pr__nfet_01v8__keta_diff_52 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_53 = {sky130_fd_pr__nfet_01v8__keta_diff_53 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_54 = {sky130_fd_pr__nfet_01v8__keta_diff_54 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_55 = {sky130_fd_pr__nfet_01v8__keta_diff_55 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_56 = {sky130_fd_pr__nfet_01v8__keta_diff_56 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_57 = {sky130_fd_pr__nfet_01v8__keta_diff_57 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_58 = {sky130_fd_pr__nfet_01v8__keta_diff_58 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_59 = {sky130_fd_pr__nfet_01v8__keta_diff_59 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_6 = {sky130_fd_pr__nfet_01v8__keta_diff_6 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_60 = {sky130_fd_pr__nfet_01v8__keta_diff_60 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_61 = {sky130_fd_pr__nfet_01v8__keta_diff_61 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_62 = {sky130_fd_pr__nfet_01v8__keta_diff_62 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_7 = {sky130_fd_pr__nfet_01v8__keta_diff_7 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_8 = {sky130_fd_pr__nfet_01v8__keta_diff_8 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__keta_diff_9 = {sky130_fd_pr__nfet_01v8__keta_diff_9 + k_nfet_keta_diff_cd*X_cd + k_nfet_keta_diff_damage*X_damage + k_nfet_keta_diff_eot*X_eot + k_nfet_keta_diff_act*X_act + k_nfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_0 = {sky130_fd_pr__nfet_01v8__kt1_diff_0 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_1 = {sky130_fd_pr__nfet_01v8__kt1_diff_1 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_10 = {sky130_fd_pr__nfet_01v8__kt1_diff_10 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_11 = {sky130_fd_pr__nfet_01v8__kt1_diff_11 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_12 = {sky130_fd_pr__nfet_01v8__kt1_diff_12 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_13 = {sky130_fd_pr__nfet_01v8__kt1_diff_13 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_14 = {sky130_fd_pr__nfet_01v8__kt1_diff_14 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_15 = {sky130_fd_pr__nfet_01v8__kt1_diff_15 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_16 = {sky130_fd_pr__nfet_01v8__kt1_diff_16 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_17 = {sky130_fd_pr__nfet_01v8__kt1_diff_17 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_18 = {sky130_fd_pr__nfet_01v8__kt1_diff_18 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_19 = {sky130_fd_pr__nfet_01v8__kt1_diff_19 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_2 = {sky130_fd_pr__nfet_01v8__kt1_diff_2 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_20 = {sky130_fd_pr__nfet_01v8__kt1_diff_20 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_21 = {sky130_fd_pr__nfet_01v8__kt1_diff_21 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_22 = {sky130_fd_pr__nfet_01v8__kt1_diff_22 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_23 = {sky130_fd_pr__nfet_01v8__kt1_diff_23 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_24 = {sky130_fd_pr__nfet_01v8__kt1_diff_24 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_25 = {sky130_fd_pr__nfet_01v8__kt1_diff_25 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_26 = {sky130_fd_pr__nfet_01v8__kt1_diff_26 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_27 = {sky130_fd_pr__nfet_01v8__kt1_diff_27 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_28 = {sky130_fd_pr__nfet_01v8__kt1_diff_28 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_29 = {sky130_fd_pr__nfet_01v8__kt1_diff_29 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_3 = {sky130_fd_pr__nfet_01v8__kt1_diff_3 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_30 = {sky130_fd_pr__nfet_01v8__kt1_diff_30 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_31 = {sky130_fd_pr__nfet_01v8__kt1_diff_31 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_32 = {sky130_fd_pr__nfet_01v8__kt1_diff_32 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_33 = {sky130_fd_pr__nfet_01v8__kt1_diff_33 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_34 = {sky130_fd_pr__nfet_01v8__kt1_diff_34 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_35 = {sky130_fd_pr__nfet_01v8__kt1_diff_35 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_36 = {sky130_fd_pr__nfet_01v8__kt1_diff_36 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_37 = {sky130_fd_pr__nfet_01v8__kt1_diff_37 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_38 = {sky130_fd_pr__nfet_01v8__kt1_diff_38 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_39 = {sky130_fd_pr__nfet_01v8__kt1_diff_39 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_4 = {sky130_fd_pr__nfet_01v8__kt1_diff_4 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_40 = {sky130_fd_pr__nfet_01v8__kt1_diff_40 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_41 = {sky130_fd_pr__nfet_01v8__kt1_diff_41 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_42 = {sky130_fd_pr__nfet_01v8__kt1_diff_42 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_43 = {sky130_fd_pr__nfet_01v8__kt1_diff_43 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_44 = {sky130_fd_pr__nfet_01v8__kt1_diff_44 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_45 = {sky130_fd_pr__nfet_01v8__kt1_diff_45 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_46 = {sky130_fd_pr__nfet_01v8__kt1_diff_46 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_47 = {sky130_fd_pr__nfet_01v8__kt1_diff_47 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_48 = {sky130_fd_pr__nfet_01v8__kt1_diff_48 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_49 = {sky130_fd_pr__nfet_01v8__kt1_diff_49 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_5 = {sky130_fd_pr__nfet_01v8__kt1_diff_5 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_50 = {sky130_fd_pr__nfet_01v8__kt1_diff_50 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_51 = {sky130_fd_pr__nfet_01v8__kt1_diff_51 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_52 = {sky130_fd_pr__nfet_01v8__kt1_diff_52 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_53 = {sky130_fd_pr__nfet_01v8__kt1_diff_53 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_54 = {sky130_fd_pr__nfet_01v8__kt1_diff_54 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_55 = {sky130_fd_pr__nfet_01v8__kt1_diff_55 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_56 = {sky130_fd_pr__nfet_01v8__kt1_diff_56 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_57 = {sky130_fd_pr__nfet_01v8__kt1_diff_57 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_58 = {sky130_fd_pr__nfet_01v8__kt1_diff_58 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_59 = {sky130_fd_pr__nfet_01v8__kt1_diff_59 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_6 = {sky130_fd_pr__nfet_01v8__kt1_diff_6 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_60 = {sky130_fd_pr__nfet_01v8__kt1_diff_60 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_61 = {sky130_fd_pr__nfet_01v8__kt1_diff_61 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_62 = {sky130_fd_pr__nfet_01v8__kt1_diff_62 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_7 = {sky130_fd_pr__nfet_01v8__kt1_diff_7 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_8 = {sky130_fd_pr__nfet_01v8__kt1_diff_8 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__kt1_diff_9 = {sky130_fd_pr__nfet_01v8__kt1_diff_9 + k_nfet_kt1_diff_cd*X_cd + k_nfet_kt1_diff_damage*X_damage + k_nfet_kt1_diff_eot*X_eot + k_nfet_kt1_diff_act*X_act + k_nfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_0 = {sky130_fd_pr__nfet_01v8__nfactor_diff_0 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_1 = {sky130_fd_pr__nfet_01v8__nfactor_diff_1 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_10 = {sky130_fd_pr__nfet_01v8__nfactor_diff_10 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_11 = {sky130_fd_pr__nfet_01v8__nfactor_diff_11 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_12 = {sky130_fd_pr__nfet_01v8__nfactor_diff_12 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_13 = {sky130_fd_pr__nfet_01v8__nfactor_diff_13 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_14 = {sky130_fd_pr__nfet_01v8__nfactor_diff_14 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_15 = {sky130_fd_pr__nfet_01v8__nfactor_diff_15 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_16 = {sky130_fd_pr__nfet_01v8__nfactor_diff_16 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_17 = {sky130_fd_pr__nfet_01v8__nfactor_diff_17 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_18 = {sky130_fd_pr__nfet_01v8__nfactor_diff_18 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_19 = {sky130_fd_pr__nfet_01v8__nfactor_diff_19 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_2 = {sky130_fd_pr__nfet_01v8__nfactor_diff_2 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_20 = {sky130_fd_pr__nfet_01v8__nfactor_diff_20 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_21 = {sky130_fd_pr__nfet_01v8__nfactor_diff_21 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_22 = {sky130_fd_pr__nfet_01v8__nfactor_diff_22 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_23 = {sky130_fd_pr__nfet_01v8__nfactor_diff_23 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_24 = {sky130_fd_pr__nfet_01v8__nfactor_diff_24 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_25 = {sky130_fd_pr__nfet_01v8__nfactor_diff_25 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_26 = {sky130_fd_pr__nfet_01v8__nfactor_diff_26 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_27 = {sky130_fd_pr__nfet_01v8__nfactor_diff_27 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_28 = {sky130_fd_pr__nfet_01v8__nfactor_diff_28 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_29 = {sky130_fd_pr__nfet_01v8__nfactor_diff_29 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_3 = {sky130_fd_pr__nfet_01v8__nfactor_diff_3 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_30 = {sky130_fd_pr__nfet_01v8__nfactor_diff_30 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_31 = {sky130_fd_pr__nfet_01v8__nfactor_diff_31 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_32 = {sky130_fd_pr__nfet_01v8__nfactor_diff_32 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_33 = {sky130_fd_pr__nfet_01v8__nfactor_diff_33 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_34 = {sky130_fd_pr__nfet_01v8__nfactor_diff_34 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_35 = {sky130_fd_pr__nfet_01v8__nfactor_diff_35 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_36 = {sky130_fd_pr__nfet_01v8__nfactor_diff_36 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_37 = {sky130_fd_pr__nfet_01v8__nfactor_diff_37 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_38 = {sky130_fd_pr__nfet_01v8__nfactor_diff_38 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_39 = {sky130_fd_pr__nfet_01v8__nfactor_diff_39 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_4 = {sky130_fd_pr__nfet_01v8__nfactor_diff_4 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_40 = {sky130_fd_pr__nfet_01v8__nfactor_diff_40 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_41 = {sky130_fd_pr__nfet_01v8__nfactor_diff_41 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_42 = {sky130_fd_pr__nfet_01v8__nfactor_diff_42 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_43 = {sky130_fd_pr__nfet_01v8__nfactor_diff_43 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_44 = {sky130_fd_pr__nfet_01v8__nfactor_diff_44 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_45 = {sky130_fd_pr__nfet_01v8__nfactor_diff_45 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_46 = {sky130_fd_pr__nfet_01v8__nfactor_diff_46 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_47 = {sky130_fd_pr__nfet_01v8__nfactor_diff_47 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_48 = {sky130_fd_pr__nfet_01v8__nfactor_diff_48 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_49 = {sky130_fd_pr__nfet_01v8__nfactor_diff_49 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_5 = {sky130_fd_pr__nfet_01v8__nfactor_diff_5 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_50 = {sky130_fd_pr__nfet_01v8__nfactor_diff_50 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_51 = {sky130_fd_pr__nfet_01v8__nfactor_diff_51 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_52 = {sky130_fd_pr__nfet_01v8__nfactor_diff_52 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_53 = {sky130_fd_pr__nfet_01v8__nfactor_diff_53 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_54 = {sky130_fd_pr__nfet_01v8__nfactor_diff_54 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_55 = {sky130_fd_pr__nfet_01v8__nfactor_diff_55 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_56 = {sky130_fd_pr__nfet_01v8__nfactor_diff_56 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_57 = {sky130_fd_pr__nfet_01v8__nfactor_diff_57 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_58 = {sky130_fd_pr__nfet_01v8__nfactor_diff_58 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_59 = {sky130_fd_pr__nfet_01v8__nfactor_diff_59 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_6 = {sky130_fd_pr__nfet_01v8__nfactor_diff_6 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_60 = {sky130_fd_pr__nfet_01v8__nfactor_diff_60 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_61 = {sky130_fd_pr__nfet_01v8__nfactor_diff_61 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_62 = {sky130_fd_pr__nfet_01v8__nfactor_diff_62 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_7 = {sky130_fd_pr__nfet_01v8__nfactor_diff_7 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_8 = {sky130_fd_pr__nfet_01v8__nfactor_diff_8 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__nfactor_diff_9 = {sky130_fd_pr__nfet_01v8__nfactor_diff_9 + k_nfet_nfactor_diff_cd*X_cd + k_nfet_nfactor_diff_damage*X_damage + k_nfet_nfactor_diff_eot*X_eot + k_nfet_nfactor_diff_act*X_act + k_nfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_0 = {sky130_fd_pr__nfet_01v8__pclm_diff_0 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_1 = {sky130_fd_pr__nfet_01v8__pclm_diff_1 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_10 = {sky130_fd_pr__nfet_01v8__pclm_diff_10 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_11 = {sky130_fd_pr__nfet_01v8__pclm_diff_11 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_12 = {sky130_fd_pr__nfet_01v8__pclm_diff_12 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_13 = {sky130_fd_pr__nfet_01v8__pclm_diff_13 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_14 = {sky130_fd_pr__nfet_01v8__pclm_diff_14 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_15 = {sky130_fd_pr__nfet_01v8__pclm_diff_15 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_16 = {sky130_fd_pr__nfet_01v8__pclm_diff_16 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_17 = {sky130_fd_pr__nfet_01v8__pclm_diff_17 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_18 = {sky130_fd_pr__nfet_01v8__pclm_diff_18 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_19 = {sky130_fd_pr__nfet_01v8__pclm_diff_19 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_2 = {sky130_fd_pr__nfet_01v8__pclm_diff_2 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_20 = {sky130_fd_pr__nfet_01v8__pclm_diff_20 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_21 = {sky130_fd_pr__nfet_01v8__pclm_diff_21 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_22 = {sky130_fd_pr__nfet_01v8__pclm_diff_22 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_23 = {sky130_fd_pr__nfet_01v8__pclm_diff_23 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_24 = {sky130_fd_pr__nfet_01v8__pclm_diff_24 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_25 = {sky130_fd_pr__nfet_01v8__pclm_diff_25 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_26 = {sky130_fd_pr__nfet_01v8__pclm_diff_26 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_27 = {sky130_fd_pr__nfet_01v8__pclm_diff_27 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_28 = {sky130_fd_pr__nfet_01v8__pclm_diff_28 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_29 = {sky130_fd_pr__nfet_01v8__pclm_diff_29 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_3 = {sky130_fd_pr__nfet_01v8__pclm_diff_3 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_30 = {sky130_fd_pr__nfet_01v8__pclm_diff_30 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_31 = {sky130_fd_pr__nfet_01v8__pclm_diff_31 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_32 = {sky130_fd_pr__nfet_01v8__pclm_diff_32 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_33 = {sky130_fd_pr__nfet_01v8__pclm_diff_33 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_34 = {sky130_fd_pr__nfet_01v8__pclm_diff_34 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_35 = {sky130_fd_pr__nfet_01v8__pclm_diff_35 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_36 = {sky130_fd_pr__nfet_01v8__pclm_diff_36 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_37 = {sky130_fd_pr__nfet_01v8__pclm_diff_37 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_38 = {sky130_fd_pr__nfet_01v8__pclm_diff_38 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_39 = {sky130_fd_pr__nfet_01v8__pclm_diff_39 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_4 = {sky130_fd_pr__nfet_01v8__pclm_diff_4 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_40 = {sky130_fd_pr__nfet_01v8__pclm_diff_40 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_41 = {sky130_fd_pr__nfet_01v8__pclm_diff_41 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_42 = {sky130_fd_pr__nfet_01v8__pclm_diff_42 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_43 = {sky130_fd_pr__nfet_01v8__pclm_diff_43 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_44 = {sky130_fd_pr__nfet_01v8__pclm_diff_44 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_45 = {sky130_fd_pr__nfet_01v8__pclm_diff_45 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_46 = {sky130_fd_pr__nfet_01v8__pclm_diff_46 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_47 = {sky130_fd_pr__nfet_01v8__pclm_diff_47 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_48 = {sky130_fd_pr__nfet_01v8__pclm_diff_48 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_49 = {sky130_fd_pr__nfet_01v8__pclm_diff_49 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_5 = {sky130_fd_pr__nfet_01v8__pclm_diff_5 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_50 = {sky130_fd_pr__nfet_01v8__pclm_diff_50 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_51 = {sky130_fd_pr__nfet_01v8__pclm_diff_51 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_52 = {sky130_fd_pr__nfet_01v8__pclm_diff_52 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_53 = {sky130_fd_pr__nfet_01v8__pclm_diff_53 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_54 = {sky130_fd_pr__nfet_01v8__pclm_diff_54 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_55 = {sky130_fd_pr__nfet_01v8__pclm_diff_55 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_56 = {sky130_fd_pr__nfet_01v8__pclm_diff_56 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_57 = {sky130_fd_pr__nfet_01v8__pclm_diff_57 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_58 = {sky130_fd_pr__nfet_01v8__pclm_diff_58 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_59 = {sky130_fd_pr__nfet_01v8__pclm_diff_59 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_6 = {sky130_fd_pr__nfet_01v8__pclm_diff_6 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_60 = {sky130_fd_pr__nfet_01v8__pclm_diff_60 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_61 = {sky130_fd_pr__nfet_01v8__pclm_diff_61 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_62 = {sky130_fd_pr__nfet_01v8__pclm_diff_62 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_7 = {sky130_fd_pr__nfet_01v8__pclm_diff_7 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_8 = {sky130_fd_pr__nfet_01v8__pclm_diff_8 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pclm_diff_9 = {sky130_fd_pr__nfet_01v8__pclm_diff_9 + k_nfet_pclm_diff_cd*X_cd + k_nfet_pclm_diff_damage*X_damage + k_nfet_pclm_diff_eot*X_eot + k_nfet_pclm_diff_act*X_act + k_nfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_0 = {sky130_fd_pr__nfet_01v8__pdits_diff_0 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_1 = {sky130_fd_pr__nfet_01v8__pdits_diff_1 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_10 = {sky130_fd_pr__nfet_01v8__pdits_diff_10 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_11 = {sky130_fd_pr__nfet_01v8__pdits_diff_11 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_12 = {sky130_fd_pr__nfet_01v8__pdits_diff_12 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_13 = {sky130_fd_pr__nfet_01v8__pdits_diff_13 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_14 = {sky130_fd_pr__nfet_01v8__pdits_diff_14 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_15 = {sky130_fd_pr__nfet_01v8__pdits_diff_15 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_16 = {sky130_fd_pr__nfet_01v8__pdits_diff_16 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_17 = {sky130_fd_pr__nfet_01v8__pdits_diff_17 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_18 = {sky130_fd_pr__nfet_01v8__pdits_diff_18 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_19 = {sky130_fd_pr__nfet_01v8__pdits_diff_19 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_2 = {sky130_fd_pr__nfet_01v8__pdits_diff_2 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_20 = {sky130_fd_pr__nfet_01v8__pdits_diff_20 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_21 = {sky130_fd_pr__nfet_01v8__pdits_diff_21 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_22 = {sky130_fd_pr__nfet_01v8__pdits_diff_22 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_23 = {sky130_fd_pr__nfet_01v8__pdits_diff_23 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_24 = {sky130_fd_pr__nfet_01v8__pdits_diff_24 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_25 = {sky130_fd_pr__nfet_01v8__pdits_diff_25 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_26 = {sky130_fd_pr__nfet_01v8__pdits_diff_26 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_27 = {sky130_fd_pr__nfet_01v8__pdits_diff_27 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_28 = {sky130_fd_pr__nfet_01v8__pdits_diff_28 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_29 = {sky130_fd_pr__nfet_01v8__pdits_diff_29 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_3 = {sky130_fd_pr__nfet_01v8__pdits_diff_3 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_30 = {sky130_fd_pr__nfet_01v8__pdits_diff_30 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_31 = {sky130_fd_pr__nfet_01v8__pdits_diff_31 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_32 = {sky130_fd_pr__nfet_01v8__pdits_diff_32 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_33 = {sky130_fd_pr__nfet_01v8__pdits_diff_33 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_34 = {sky130_fd_pr__nfet_01v8__pdits_diff_34 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_35 = {sky130_fd_pr__nfet_01v8__pdits_diff_35 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_36 = {sky130_fd_pr__nfet_01v8__pdits_diff_36 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_37 = {sky130_fd_pr__nfet_01v8__pdits_diff_37 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_38 = {sky130_fd_pr__nfet_01v8__pdits_diff_38 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_39 = {sky130_fd_pr__nfet_01v8__pdits_diff_39 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_4 = {sky130_fd_pr__nfet_01v8__pdits_diff_4 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_40 = {sky130_fd_pr__nfet_01v8__pdits_diff_40 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_41 = {sky130_fd_pr__nfet_01v8__pdits_diff_41 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_42 = {sky130_fd_pr__nfet_01v8__pdits_diff_42 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_43 = {sky130_fd_pr__nfet_01v8__pdits_diff_43 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_44 = {sky130_fd_pr__nfet_01v8__pdits_diff_44 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_45 = {sky130_fd_pr__nfet_01v8__pdits_diff_45 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_46 = {sky130_fd_pr__nfet_01v8__pdits_diff_46 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_47 = {sky130_fd_pr__nfet_01v8__pdits_diff_47 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_48 = {sky130_fd_pr__nfet_01v8__pdits_diff_48 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_49 = {sky130_fd_pr__nfet_01v8__pdits_diff_49 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_5 = {sky130_fd_pr__nfet_01v8__pdits_diff_5 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_50 = {sky130_fd_pr__nfet_01v8__pdits_diff_50 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_51 = {sky130_fd_pr__nfet_01v8__pdits_diff_51 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_52 = {sky130_fd_pr__nfet_01v8__pdits_diff_52 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_53 = {sky130_fd_pr__nfet_01v8__pdits_diff_53 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_54 = {sky130_fd_pr__nfet_01v8__pdits_diff_54 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_55 = {sky130_fd_pr__nfet_01v8__pdits_diff_55 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_56 = {sky130_fd_pr__nfet_01v8__pdits_diff_56 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_57 = {sky130_fd_pr__nfet_01v8__pdits_diff_57 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_58 = {sky130_fd_pr__nfet_01v8__pdits_diff_58 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_59 = {sky130_fd_pr__nfet_01v8__pdits_diff_59 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_6 = {sky130_fd_pr__nfet_01v8__pdits_diff_6 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_60 = {sky130_fd_pr__nfet_01v8__pdits_diff_60 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_61 = {sky130_fd_pr__nfet_01v8__pdits_diff_61 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_62 = {sky130_fd_pr__nfet_01v8__pdits_diff_62 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_7 = {sky130_fd_pr__nfet_01v8__pdits_diff_7 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_8 = {sky130_fd_pr__nfet_01v8__pdits_diff_8 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pdits_diff_9 = {sky130_fd_pr__nfet_01v8__pdits_diff_9 + k_nfet_pdits_diff_cd*X_cd + k_nfet_pdits_diff_damage*X_damage + k_nfet_pdits_diff_eot*X_eot + k_nfet_pdits_diff_act*X_act + k_nfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_0 = {sky130_fd_pr__nfet_01v8__pditsd_diff_0 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_1 = {sky130_fd_pr__nfet_01v8__pditsd_diff_1 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_10 = {sky130_fd_pr__nfet_01v8__pditsd_diff_10 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_11 = {sky130_fd_pr__nfet_01v8__pditsd_diff_11 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_12 = {sky130_fd_pr__nfet_01v8__pditsd_diff_12 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_13 = {sky130_fd_pr__nfet_01v8__pditsd_diff_13 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_14 = {sky130_fd_pr__nfet_01v8__pditsd_diff_14 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_15 = {sky130_fd_pr__nfet_01v8__pditsd_diff_15 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_16 = {sky130_fd_pr__nfet_01v8__pditsd_diff_16 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_17 = {sky130_fd_pr__nfet_01v8__pditsd_diff_17 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_18 = {sky130_fd_pr__nfet_01v8__pditsd_diff_18 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_19 = {sky130_fd_pr__nfet_01v8__pditsd_diff_19 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_2 = {sky130_fd_pr__nfet_01v8__pditsd_diff_2 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_20 = {sky130_fd_pr__nfet_01v8__pditsd_diff_20 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_21 = {sky130_fd_pr__nfet_01v8__pditsd_diff_21 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_22 = {sky130_fd_pr__nfet_01v8__pditsd_diff_22 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_23 = {sky130_fd_pr__nfet_01v8__pditsd_diff_23 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_24 = {sky130_fd_pr__nfet_01v8__pditsd_diff_24 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_25 = {sky130_fd_pr__nfet_01v8__pditsd_diff_25 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_26 = {sky130_fd_pr__nfet_01v8__pditsd_diff_26 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_27 = {sky130_fd_pr__nfet_01v8__pditsd_diff_27 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_28 = {sky130_fd_pr__nfet_01v8__pditsd_diff_28 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_29 = {sky130_fd_pr__nfet_01v8__pditsd_diff_29 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_3 = {sky130_fd_pr__nfet_01v8__pditsd_diff_3 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_30 = {sky130_fd_pr__nfet_01v8__pditsd_diff_30 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_31 = {sky130_fd_pr__nfet_01v8__pditsd_diff_31 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_32 = {sky130_fd_pr__nfet_01v8__pditsd_diff_32 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_33 = {sky130_fd_pr__nfet_01v8__pditsd_diff_33 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_34 = {sky130_fd_pr__nfet_01v8__pditsd_diff_34 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_35 = {sky130_fd_pr__nfet_01v8__pditsd_diff_35 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_36 = {sky130_fd_pr__nfet_01v8__pditsd_diff_36 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_37 = {sky130_fd_pr__nfet_01v8__pditsd_diff_37 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_38 = {sky130_fd_pr__nfet_01v8__pditsd_diff_38 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_39 = {sky130_fd_pr__nfet_01v8__pditsd_diff_39 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_4 = {sky130_fd_pr__nfet_01v8__pditsd_diff_4 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_40 = {sky130_fd_pr__nfet_01v8__pditsd_diff_40 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_41 = {sky130_fd_pr__nfet_01v8__pditsd_diff_41 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_42 = {sky130_fd_pr__nfet_01v8__pditsd_diff_42 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_43 = {sky130_fd_pr__nfet_01v8__pditsd_diff_43 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_44 = {sky130_fd_pr__nfet_01v8__pditsd_diff_44 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_45 = {sky130_fd_pr__nfet_01v8__pditsd_diff_45 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_46 = {sky130_fd_pr__nfet_01v8__pditsd_diff_46 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_47 = {sky130_fd_pr__nfet_01v8__pditsd_diff_47 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_48 = {sky130_fd_pr__nfet_01v8__pditsd_diff_48 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_49 = {sky130_fd_pr__nfet_01v8__pditsd_diff_49 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_5 = {sky130_fd_pr__nfet_01v8__pditsd_diff_5 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_50 = {sky130_fd_pr__nfet_01v8__pditsd_diff_50 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_51 = {sky130_fd_pr__nfet_01v8__pditsd_diff_51 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_52 = {sky130_fd_pr__nfet_01v8__pditsd_diff_52 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_53 = {sky130_fd_pr__nfet_01v8__pditsd_diff_53 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_54 = {sky130_fd_pr__nfet_01v8__pditsd_diff_54 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_55 = {sky130_fd_pr__nfet_01v8__pditsd_diff_55 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_56 = {sky130_fd_pr__nfet_01v8__pditsd_diff_56 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_57 = {sky130_fd_pr__nfet_01v8__pditsd_diff_57 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_58 = {sky130_fd_pr__nfet_01v8__pditsd_diff_58 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_59 = {sky130_fd_pr__nfet_01v8__pditsd_diff_59 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_6 = {sky130_fd_pr__nfet_01v8__pditsd_diff_6 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_60 = {sky130_fd_pr__nfet_01v8__pditsd_diff_60 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_61 = {sky130_fd_pr__nfet_01v8__pditsd_diff_61 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_62 = {sky130_fd_pr__nfet_01v8__pditsd_diff_62 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_7 = {sky130_fd_pr__nfet_01v8__pditsd_diff_7 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_8 = {sky130_fd_pr__nfet_01v8__pditsd_diff_8 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__pditsd_diff_9 = {sky130_fd_pr__nfet_01v8__pditsd_diff_9 + k_nfet_pditsd_diff_cd*X_cd + k_nfet_pditsd_diff_damage*X_damage + k_nfet_pditsd_diff_eot*X_eot + k_nfet_pditsd_diff_act*X_act + k_nfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_0 = {sky130_fd_pr__nfet_01v8__rdsw_diff_0 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_1 = {sky130_fd_pr__nfet_01v8__rdsw_diff_1 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_10 = {sky130_fd_pr__nfet_01v8__rdsw_diff_10 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_11 = {sky130_fd_pr__nfet_01v8__rdsw_diff_11 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_12 = {sky130_fd_pr__nfet_01v8__rdsw_diff_12 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_13 = {sky130_fd_pr__nfet_01v8__rdsw_diff_13 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_14 = {sky130_fd_pr__nfet_01v8__rdsw_diff_14 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_15 = {sky130_fd_pr__nfet_01v8__rdsw_diff_15 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_16 = {sky130_fd_pr__nfet_01v8__rdsw_diff_16 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_17 = {sky130_fd_pr__nfet_01v8__rdsw_diff_17 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_18 = {sky130_fd_pr__nfet_01v8__rdsw_diff_18 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_19 = {sky130_fd_pr__nfet_01v8__rdsw_diff_19 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_2 = {sky130_fd_pr__nfet_01v8__rdsw_diff_2 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_20 = {sky130_fd_pr__nfet_01v8__rdsw_diff_20 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_21 = {sky130_fd_pr__nfet_01v8__rdsw_diff_21 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_22 = {sky130_fd_pr__nfet_01v8__rdsw_diff_22 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_23 = {sky130_fd_pr__nfet_01v8__rdsw_diff_23 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_24 = {sky130_fd_pr__nfet_01v8__rdsw_diff_24 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_25 = {sky130_fd_pr__nfet_01v8__rdsw_diff_25 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_26 = {sky130_fd_pr__nfet_01v8__rdsw_diff_26 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_27 = {sky130_fd_pr__nfet_01v8__rdsw_diff_27 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_28 = {sky130_fd_pr__nfet_01v8__rdsw_diff_28 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_29 = {sky130_fd_pr__nfet_01v8__rdsw_diff_29 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_3 = {sky130_fd_pr__nfet_01v8__rdsw_diff_3 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_30 = {sky130_fd_pr__nfet_01v8__rdsw_diff_30 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_31 = {sky130_fd_pr__nfet_01v8__rdsw_diff_31 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_32 = {sky130_fd_pr__nfet_01v8__rdsw_diff_32 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_33 = {sky130_fd_pr__nfet_01v8__rdsw_diff_33 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_34 = {sky130_fd_pr__nfet_01v8__rdsw_diff_34 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_35 = {sky130_fd_pr__nfet_01v8__rdsw_diff_35 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_36 = {sky130_fd_pr__nfet_01v8__rdsw_diff_36 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_37 = {sky130_fd_pr__nfet_01v8__rdsw_diff_37 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_38 = {sky130_fd_pr__nfet_01v8__rdsw_diff_38 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_39 = {sky130_fd_pr__nfet_01v8__rdsw_diff_39 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_4 = {sky130_fd_pr__nfet_01v8__rdsw_diff_4 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_40 = {sky130_fd_pr__nfet_01v8__rdsw_diff_40 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_41 = {sky130_fd_pr__nfet_01v8__rdsw_diff_41 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_42 = {sky130_fd_pr__nfet_01v8__rdsw_diff_42 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_43 = {sky130_fd_pr__nfet_01v8__rdsw_diff_43 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_44 = {sky130_fd_pr__nfet_01v8__rdsw_diff_44 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_45 = {sky130_fd_pr__nfet_01v8__rdsw_diff_45 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_46 = {sky130_fd_pr__nfet_01v8__rdsw_diff_46 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_47 = {sky130_fd_pr__nfet_01v8__rdsw_diff_47 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_48 = {sky130_fd_pr__nfet_01v8__rdsw_diff_48 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_49 = {sky130_fd_pr__nfet_01v8__rdsw_diff_49 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_5 = {sky130_fd_pr__nfet_01v8__rdsw_diff_5 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_50 = {sky130_fd_pr__nfet_01v8__rdsw_diff_50 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_51 = {sky130_fd_pr__nfet_01v8__rdsw_diff_51 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_52 = {sky130_fd_pr__nfet_01v8__rdsw_diff_52 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_53 = {sky130_fd_pr__nfet_01v8__rdsw_diff_53 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_54 = {sky130_fd_pr__nfet_01v8__rdsw_diff_54 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_55 = {sky130_fd_pr__nfet_01v8__rdsw_diff_55 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_56 = {sky130_fd_pr__nfet_01v8__rdsw_diff_56 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_57 = {sky130_fd_pr__nfet_01v8__rdsw_diff_57 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_58 = {sky130_fd_pr__nfet_01v8__rdsw_diff_58 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_59 = {sky130_fd_pr__nfet_01v8__rdsw_diff_59 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_6 = {sky130_fd_pr__nfet_01v8__rdsw_diff_6 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_60 = {sky130_fd_pr__nfet_01v8__rdsw_diff_60 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_61 = {sky130_fd_pr__nfet_01v8__rdsw_diff_61 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_62 = {sky130_fd_pr__nfet_01v8__rdsw_diff_62 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_7 = {sky130_fd_pr__nfet_01v8__rdsw_diff_7 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_8 = {sky130_fd_pr__nfet_01v8__rdsw_diff_8 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__rdsw_diff_9 = {sky130_fd_pr__nfet_01v8__rdsw_diff_9 + k_nfet_rdsw_diff_cd*X_cd + k_nfet_rdsw_diff_damage*X_damage + k_nfet_rdsw_diff_eot*X_eot + k_nfet_rdsw_diff_act*X_act + k_nfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_0 = {sky130_fd_pr__nfet_01v8__tvoff_diff_0 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_1 = {sky130_fd_pr__nfet_01v8__tvoff_diff_1 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_10 = {sky130_fd_pr__nfet_01v8__tvoff_diff_10 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_11 = {sky130_fd_pr__nfet_01v8__tvoff_diff_11 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_12 = {sky130_fd_pr__nfet_01v8__tvoff_diff_12 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_13 = {sky130_fd_pr__nfet_01v8__tvoff_diff_13 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_14 = {sky130_fd_pr__nfet_01v8__tvoff_diff_14 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_15 = {sky130_fd_pr__nfet_01v8__tvoff_diff_15 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_16 = {sky130_fd_pr__nfet_01v8__tvoff_diff_16 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_17 = {sky130_fd_pr__nfet_01v8__tvoff_diff_17 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_18 = {sky130_fd_pr__nfet_01v8__tvoff_diff_18 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_19 = {sky130_fd_pr__nfet_01v8__tvoff_diff_19 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_2 = {sky130_fd_pr__nfet_01v8__tvoff_diff_2 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_20 = {sky130_fd_pr__nfet_01v8__tvoff_diff_20 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_21 = {sky130_fd_pr__nfet_01v8__tvoff_diff_21 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_22 = {sky130_fd_pr__nfet_01v8__tvoff_diff_22 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_23 = {sky130_fd_pr__nfet_01v8__tvoff_diff_23 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_24 = {sky130_fd_pr__nfet_01v8__tvoff_diff_24 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_25 = {sky130_fd_pr__nfet_01v8__tvoff_diff_25 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_26 = {sky130_fd_pr__nfet_01v8__tvoff_diff_26 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_27 = {sky130_fd_pr__nfet_01v8__tvoff_diff_27 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_28 = {sky130_fd_pr__nfet_01v8__tvoff_diff_28 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_29 = {sky130_fd_pr__nfet_01v8__tvoff_diff_29 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_3 = {sky130_fd_pr__nfet_01v8__tvoff_diff_3 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_30 = {sky130_fd_pr__nfet_01v8__tvoff_diff_30 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_31 = {sky130_fd_pr__nfet_01v8__tvoff_diff_31 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_32 = {sky130_fd_pr__nfet_01v8__tvoff_diff_32 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_33 = {sky130_fd_pr__nfet_01v8__tvoff_diff_33 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_34 = {sky130_fd_pr__nfet_01v8__tvoff_diff_34 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_35 = {sky130_fd_pr__nfet_01v8__tvoff_diff_35 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_36 = {sky130_fd_pr__nfet_01v8__tvoff_diff_36 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_37 = {sky130_fd_pr__nfet_01v8__tvoff_diff_37 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_38 = {sky130_fd_pr__nfet_01v8__tvoff_diff_38 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_39 = {sky130_fd_pr__nfet_01v8__tvoff_diff_39 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_4 = {sky130_fd_pr__nfet_01v8__tvoff_diff_4 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_40 = {sky130_fd_pr__nfet_01v8__tvoff_diff_40 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_41 = {sky130_fd_pr__nfet_01v8__tvoff_diff_41 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_42 = {sky130_fd_pr__nfet_01v8__tvoff_diff_42 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_43 = {sky130_fd_pr__nfet_01v8__tvoff_diff_43 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_44 = {sky130_fd_pr__nfet_01v8__tvoff_diff_44 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_45 = {sky130_fd_pr__nfet_01v8__tvoff_diff_45 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_46 = {sky130_fd_pr__nfet_01v8__tvoff_diff_46 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_47 = {sky130_fd_pr__nfet_01v8__tvoff_diff_47 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_48 = {sky130_fd_pr__nfet_01v8__tvoff_diff_48 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_49 = {sky130_fd_pr__nfet_01v8__tvoff_diff_49 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_5 = {sky130_fd_pr__nfet_01v8__tvoff_diff_5 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_50 = {sky130_fd_pr__nfet_01v8__tvoff_diff_50 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_51 = {sky130_fd_pr__nfet_01v8__tvoff_diff_51 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_52 = {sky130_fd_pr__nfet_01v8__tvoff_diff_52 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_53 = {sky130_fd_pr__nfet_01v8__tvoff_diff_53 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_54 = {sky130_fd_pr__nfet_01v8__tvoff_diff_54 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_55 = {sky130_fd_pr__nfet_01v8__tvoff_diff_55 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_56 = {sky130_fd_pr__nfet_01v8__tvoff_diff_56 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_57 = {sky130_fd_pr__nfet_01v8__tvoff_diff_57 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_58 = {sky130_fd_pr__nfet_01v8__tvoff_diff_58 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_59 = {sky130_fd_pr__nfet_01v8__tvoff_diff_59 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_6 = {sky130_fd_pr__nfet_01v8__tvoff_diff_6 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_60 = {sky130_fd_pr__nfet_01v8__tvoff_diff_60 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_61 = {sky130_fd_pr__nfet_01v8__tvoff_diff_61 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_62 = {sky130_fd_pr__nfet_01v8__tvoff_diff_62 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_7 = {sky130_fd_pr__nfet_01v8__tvoff_diff_7 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_8 = {sky130_fd_pr__nfet_01v8__tvoff_diff_8 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__tvoff_diff_9 = {sky130_fd_pr__nfet_01v8__tvoff_diff_9 + k_nfet_tvoff_diff_cd*X_cd + k_nfet_tvoff_diff_damage*X_damage + k_nfet_tvoff_diff_eot*X_eot + k_nfet_tvoff_diff_act*X_act + k_nfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_0 = {sky130_fd_pr__nfet_01v8__u0_diff_0 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_1 = {sky130_fd_pr__nfet_01v8__u0_diff_1 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_10 = {sky130_fd_pr__nfet_01v8__u0_diff_10 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_11 = {sky130_fd_pr__nfet_01v8__u0_diff_11 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_12 = {sky130_fd_pr__nfet_01v8__u0_diff_12 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_13 = {sky130_fd_pr__nfet_01v8__u0_diff_13 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_14 = {sky130_fd_pr__nfet_01v8__u0_diff_14 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_15 = {sky130_fd_pr__nfet_01v8__u0_diff_15 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_16 = {sky130_fd_pr__nfet_01v8__u0_diff_16 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_17 = {sky130_fd_pr__nfet_01v8__u0_diff_17 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_18 = {sky130_fd_pr__nfet_01v8__u0_diff_18 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_19 = {sky130_fd_pr__nfet_01v8__u0_diff_19 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_2 = {sky130_fd_pr__nfet_01v8__u0_diff_2 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_20 = {sky130_fd_pr__nfet_01v8__u0_diff_20 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_21 = {sky130_fd_pr__nfet_01v8__u0_diff_21 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_22 = {sky130_fd_pr__nfet_01v8__u0_diff_22 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_23 = {sky130_fd_pr__nfet_01v8__u0_diff_23 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_24 = {sky130_fd_pr__nfet_01v8__u0_diff_24 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_25 = {sky130_fd_pr__nfet_01v8__u0_diff_25 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_26 = {sky130_fd_pr__nfet_01v8__u0_diff_26 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_27 = {sky130_fd_pr__nfet_01v8__u0_diff_27 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_28 = {sky130_fd_pr__nfet_01v8__u0_diff_28 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_29 = {sky130_fd_pr__nfet_01v8__u0_diff_29 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_3 = {sky130_fd_pr__nfet_01v8__u0_diff_3 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_30 = {sky130_fd_pr__nfet_01v8__u0_diff_30 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_31 = {sky130_fd_pr__nfet_01v8__u0_diff_31 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_32 = {sky130_fd_pr__nfet_01v8__u0_diff_32 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_33 = {sky130_fd_pr__nfet_01v8__u0_diff_33 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_34 = {sky130_fd_pr__nfet_01v8__u0_diff_34 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_35 = {sky130_fd_pr__nfet_01v8__u0_diff_35 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_36 = {sky130_fd_pr__nfet_01v8__u0_diff_36 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_37 = {sky130_fd_pr__nfet_01v8__u0_diff_37 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_38 = {sky130_fd_pr__nfet_01v8__u0_diff_38 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_39 = {sky130_fd_pr__nfet_01v8__u0_diff_39 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_4 = {sky130_fd_pr__nfet_01v8__u0_diff_4 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_40 = {sky130_fd_pr__nfet_01v8__u0_diff_40 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_41 = {sky130_fd_pr__nfet_01v8__u0_diff_41 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_42 = {sky130_fd_pr__nfet_01v8__u0_diff_42 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_43 = {sky130_fd_pr__nfet_01v8__u0_diff_43 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_44 = {sky130_fd_pr__nfet_01v8__u0_diff_44 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_45 = {sky130_fd_pr__nfet_01v8__u0_diff_45 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_46 = {sky130_fd_pr__nfet_01v8__u0_diff_46 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_47 = {sky130_fd_pr__nfet_01v8__u0_diff_47 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_48 = {sky130_fd_pr__nfet_01v8__u0_diff_48 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_49 = {sky130_fd_pr__nfet_01v8__u0_diff_49 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_5 = {sky130_fd_pr__nfet_01v8__u0_diff_5 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_50 = {sky130_fd_pr__nfet_01v8__u0_diff_50 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_51 = {sky130_fd_pr__nfet_01v8__u0_diff_51 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_52 = {sky130_fd_pr__nfet_01v8__u0_diff_52 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_53 = {sky130_fd_pr__nfet_01v8__u0_diff_53 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_54 = {sky130_fd_pr__nfet_01v8__u0_diff_54 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_55 = {sky130_fd_pr__nfet_01v8__u0_diff_55 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_56 = {sky130_fd_pr__nfet_01v8__u0_diff_56 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_57 = {sky130_fd_pr__nfet_01v8__u0_diff_57 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_58 = {sky130_fd_pr__nfet_01v8__u0_diff_58 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_59 = {sky130_fd_pr__nfet_01v8__u0_diff_59 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_6 = {sky130_fd_pr__nfet_01v8__u0_diff_6 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_60 = {sky130_fd_pr__nfet_01v8__u0_diff_60 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_61 = {sky130_fd_pr__nfet_01v8__u0_diff_61 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_62 = {sky130_fd_pr__nfet_01v8__u0_diff_62 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_7 = {sky130_fd_pr__nfet_01v8__u0_diff_7 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_8 = {sky130_fd_pr__nfet_01v8__u0_diff_8 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__u0_diff_9 = {sky130_fd_pr__nfet_01v8__u0_diff_9 + k_nfet_u0_diff_cd*X_cd + k_nfet_u0_diff_damage*X_damage + k_nfet_u0_diff_eot*X_eot + k_nfet_u0_diff_act*X_act + k_nfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_0 = {sky130_fd_pr__nfet_01v8__ua_diff_0 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_1 = {sky130_fd_pr__nfet_01v8__ua_diff_1 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_10 = {sky130_fd_pr__nfet_01v8__ua_diff_10 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_11 = {sky130_fd_pr__nfet_01v8__ua_diff_11 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_12 = {sky130_fd_pr__nfet_01v8__ua_diff_12 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_13 = {sky130_fd_pr__nfet_01v8__ua_diff_13 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_14 = {sky130_fd_pr__nfet_01v8__ua_diff_14 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_15 = {sky130_fd_pr__nfet_01v8__ua_diff_15 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_16 = {sky130_fd_pr__nfet_01v8__ua_diff_16 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_17 = {sky130_fd_pr__nfet_01v8__ua_diff_17 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_18 = {sky130_fd_pr__nfet_01v8__ua_diff_18 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_19 = {sky130_fd_pr__nfet_01v8__ua_diff_19 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_2 = {sky130_fd_pr__nfet_01v8__ua_diff_2 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_20 = {sky130_fd_pr__nfet_01v8__ua_diff_20 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_21 = {sky130_fd_pr__nfet_01v8__ua_diff_21 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_22 = {sky130_fd_pr__nfet_01v8__ua_diff_22 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_23 = {sky130_fd_pr__nfet_01v8__ua_diff_23 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_24 = {sky130_fd_pr__nfet_01v8__ua_diff_24 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_25 = {sky130_fd_pr__nfet_01v8__ua_diff_25 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_26 = {sky130_fd_pr__nfet_01v8__ua_diff_26 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_27 = {sky130_fd_pr__nfet_01v8__ua_diff_27 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_28 = {sky130_fd_pr__nfet_01v8__ua_diff_28 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_29 = {sky130_fd_pr__nfet_01v8__ua_diff_29 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_3 = {sky130_fd_pr__nfet_01v8__ua_diff_3 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_30 = {sky130_fd_pr__nfet_01v8__ua_diff_30 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_31 = {sky130_fd_pr__nfet_01v8__ua_diff_31 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_32 = {sky130_fd_pr__nfet_01v8__ua_diff_32 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_33 = {sky130_fd_pr__nfet_01v8__ua_diff_33 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_34 = {sky130_fd_pr__nfet_01v8__ua_diff_34 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_35 = {sky130_fd_pr__nfet_01v8__ua_diff_35 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_36 = {sky130_fd_pr__nfet_01v8__ua_diff_36 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_37 = {sky130_fd_pr__nfet_01v8__ua_diff_37 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_38 = {sky130_fd_pr__nfet_01v8__ua_diff_38 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_39 = {sky130_fd_pr__nfet_01v8__ua_diff_39 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_4 = {sky130_fd_pr__nfet_01v8__ua_diff_4 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_40 = {sky130_fd_pr__nfet_01v8__ua_diff_40 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_41 = {sky130_fd_pr__nfet_01v8__ua_diff_41 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_42 = {sky130_fd_pr__nfet_01v8__ua_diff_42 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_43 = {sky130_fd_pr__nfet_01v8__ua_diff_43 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_44 = {sky130_fd_pr__nfet_01v8__ua_diff_44 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_45 = {sky130_fd_pr__nfet_01v8__ua_diff_45 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_46 = {sky130_fd_pr__nfet_01v8__ua_diff_46 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_47 = {sky130_fd_pr__nfet_01v8__ua_diff_47 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_48 = {sky130_fd_pr__nfet_01v8__ua_diff_48 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_49 = {sky130_fd_pr__nfet_01v8__ua_diff_49 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_5 = {sky130_fd_pr__nfet_01v8__ua_diff_5 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_50 = {sky130_fd_pr__nfet_01v8__ua_diff_50 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_51 = {sky130_fd_pr__nfet_01v8__ua_diff_51 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_52 = {sky130_fd_pr__nfet_01v8__ua_diff_52 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_53 = {sky130_fd_pr__nfet_01v8__ua_diff_53 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_54 = {sky130_fd_pr__nfet_01v8__ua_diff_54 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_55 = {sky130_fd_pr__nfet_01v8__ua_diff_55 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_56 = {sky130_fd_pr__nfet_01v8__ua_diff_56 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_57 = {sky130_fd_pr__nfet_01v8__ua_diff_57 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_58 = {sky130_fd_pr__nfet_01v8__ua_diff_58 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_59 = {sky130_fd_pr__nfet_01v8__ua_diff_59 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_6 = {sky130_fd_pr__nfet_01v8__ua_diff_6 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_60 = {sky130_fd_pr__nfet_01v8__ua_diff_60 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_61 = {sky130_fd_pr__nfet_01v8__ua_diff_61 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_62 = {sky130_fd_pr__nfet_01v8__ua_diff_62 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_7 = {sky130_fd_pr__nfet_01v8__ua_diff_7 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_8 = {sky130_fd_pr__nfet_01v8__ua_diff_8 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ua_diff_9 = {sky130_fd_pr__nfet_01v8__ua_diff_9 + k_nfet_ua_diff_cd*X_cd + k_nfet_ua_diff_damage*X_damage + k_nfet_ua_diff_eot*X_eot + k_nfet_ua_diff_act*X_act + k_nfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_0 = {sky130_fd_pr__nfet_01v8__ub_diff_0 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_1 = {sky130_fd_pr__nfet_01v8__ub_diff_1 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_10 = {sky130_fd_pr__nfet_01v8__ub_diff_10 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_11 = {sky130_fd_pr__nfet_01v8__ub_diff_11 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_12 = {sky130_fd_pr__nfet_01v8__ub_diff_12 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_13 = {sky130_fd_pr__nfet_01v8__ub_diff_13 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_14 = {sky130_fd_pr__nfet_01v8__ub_diff_14 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_15 = {sky130_fd_pr__nfet_01v8__ub_diff_15 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_16 = {sky130_fd_pr__nfet_01v8__ub_diff_16 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_17 = {sky130_fd_pr__nfet_01v8__ub_diff_17 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_18 = {sky130_fd_pr__nfet_01v8__ub_diff_18 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_19 = {sky130_fd_pr__nfet_01v8__ub_diff_19 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_2 = {sky130_fd_pr__nfet_01v8__ub_diff_2 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_20 = {sky130_fd_pr__nfet_01v8__ub_diff_20 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_21 = {sky130_fd_pr__nfet_01v8__ub_diff_21 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_22 = {sky130_fd_pr__nfet_01v8__ub_diff_22 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_23 = {sky130_fd_pr__nfet_01v8__ub_diff_23 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_24 = {sky130_fd_pr__nfet_01v8__ub_diff_24 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_25 = {sky130_fd_pr__nfet_01v8__ub_diff_25 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_26 = {sky130_fd_pr__nfet_01v8__ub_diff_26 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_27 = {sky130_fd_pr__nfet_01v8__ub_diff_27 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_28 = {sky130_fd_pr__nfet_01v8__ub_diff_28 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_29 = {sky130_fd_pr__nfet_01v8__ub_diff_29 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_3 = {sky130_fd_pr__nfet_01v8__ub_diff_3 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_30 = {sky130_fd_pr__nfet_01v8__ub_diff_30 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_31 = {sky130_fd_pr__nfet_01v8__ub_diff_31 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_32 = {sky130_fd_pr__nfet_01v8__ub_diff_32 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_33 = {sky130_fd_pr__nfet_01v8__ub_diff_33 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_34 = {sky130_fd_pr__nfet_01v8__ub_diff_34 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_35 = {sky130_fd_pr__nfet_01v8__ub_diff_35 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_36 = {sky130_fd_pr__nfet_01v8__ub_diff_36 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_37 = {sky130_fd_pr__nfet_01v8__ub_diff_37 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_38 = {sky130_fd_pr__nfet_01v8__ub_diff_38 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_39 = {sky130_fd_pr__nfet_01v8__ub_diff_39 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_4 = {sky130_fd_pr__nfet_01v8__ub_diff_4 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_40 = {sky130_fd_pr__nfet_01v8__ub_diff_40 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_41 = {sky130_fd_pr__nfet_01v8__ub_diff_41 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_42 = {sky130_fd_pr__nfet_01v8__ub_diff_42 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_43 = {sky130_fd_pr__nfet_01v8__ub_diff_43 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_44 = {sky130_fd_pr__nfet_01v8__ub_diff_44 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_45 = {sky130_fd_pr__nfet_01v8__ub_diff_45 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_46 = {sky130_fd_pr__nfet_01v8__ub_diff_46 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_47 = {sky130_fd_pr__nfet_01v8__ub_diff_47 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_48 = {sky130_fd_pr__nfet_01v8__ub_diff_48 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_49 = {sky130_fd_pr__nfet_01v8__ub_diff_49 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_5 = {sky130_fd_pr__nfet_01v8__ub_diff_5 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_50 = {sky130_fd_pr__nfet_01v8__ub_diff_50 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_51 = {sky130_fd_pr__nfet_01v8__ub_diff_51 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_52 = {sky130_fd_pr__nfet_01v8__ub_diff_52 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_53 = {sky130_fd_pr__nfet_01v8__ub_diff_53 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_54 = {sky130_fd_pr__nfet_01v8__ub_diff_54 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_55 = {sky130_fd_pr__nfet_01v8__ub_diff_55 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_56 = {sky130_fd_pr__nfet_01v8__ub_diff_56 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_57 = {sky130_fd_pr__nfet_01v8__ub_diff_57 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_58 = {sky130_fd_pr__nfet_01v8__ub_diff_58 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_59 = {sky130_fd_pr__nfet_01v8__ub_diff_59 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_6 = {sky130_fd_pr__nfet_01v8__ub_diff_6 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_60 = {sky130_fd_pr__nfet_01v8__ub_diff_60 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_61 = {sky130_fd_pr__nfet_01v8__ub_diff_61 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_62 = {sky130_fd_pr__nfet_01v8__ub_diff_62 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_7 = {sky130_fd_pr__nfet_01v8__ub_diff_7 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_8 = {sky130_fd_pr__nfet_01v8__ub_diff_8 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__ub_diff_9 = {sky130_fd_pr__nfet_01v8__ub_diff_9 + k_nfet_ub_diff_cd*X_cd + k_nfet_ub_diff_damage*X_damage + k_nfet_ub_diff_eot*X_eot + k_nfet_ub_diff_act*X_act + k_nfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_0 = {sky130_fd_pr__nfet_01v8__voff_diff_0 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_1 = {sky130_fd_pr__nfet_01v8__voff_diff_1 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_10 = {sky130_fd_pr__nfet_01v8__voff_diff_10 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_11 = {sky130_fd_pr__nfet_01v8__voff_diff_11 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_12 = {sky130_fd_pr__nfet_01v8__voff_diff_12 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_13 = {sky130_fd_pr__nfet_01v8__voff_diff_13 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_14 = {sky130_fd_pr__nfet_01v8__voff_diff_14 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_15 = {sky130_fd_pr__nfet_01v8__voff_diff_15 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_16 = {sky130_fd_pr__nfet_01v8__voff_diff_16 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_17 = {sky130_fd_pr__nfet_01v8__voff_diff_17 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_18 = {sky130_fd_pr__nfet_01v8__voff_diff_18 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_19 = {sky130_fd_pr__nfet_01v8__voff_diff_19 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_2 = {sky130_fd_pr__nfet_01v8__voff_diff_2 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_20 = {sky130_fd_pr__nfet_01v8__voff_diff_20 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_21 = {sky130_fd_pr__nfet_01v8__voff_diff_21 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_22 = {sky130_fd_pr__nfet_01v8__voff_diff_22 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_23 = {sky130_fd_pr__nfet_01v8__voff_diff_23 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_24 = {sky130_fd_pr__nfet_01v8__voff_diff_24 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_25 = {sky130_fd_pr__nfet_01v8__voff_diff_25 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_26 = {sky130_fd_pr__nfet_01v8__voff_diff_26 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_27 = {sky130_fd_pr__nfet_01v8__voff_diff_27 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_28 = {sky130_fd_pr__nfet_01v8__voff_diff_28 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_29 = {sky130_fd_pr__nfet_01v8__voff_diff_29 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_3 = {sky130_fd_pr__nfet_01v8__voff_diff_3 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_30 = {sky130_fd_pr__nfet_01v8__voff_diff_30 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_31 = {sky130_fd_pr__nfet_01v8__voff_diff_31 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_32 = {sky130_fd_pr__nfet_01v8__voff_diff_32 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_33 = {sky130_fd_pr__nfet_01v8__voff_diff_33 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_34 = {sky130_fd_pr__nfet_01v8__voff_diff_34 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_35 = {sky130_fd_pr__nfet_01v8__voff_diff_35 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_36 = {sky130_fd_pr__nfet_01v8__voff_diff_36 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_37 = {sky130_fd_pr__nfet_01v8__voff_diff_37 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_38 = {sky130_fd_pr__nfet_01v8__voff_diff_38 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_39 = {sky130_fd_pr__nfet_01v8__voff_diff_39 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_4 = {sky130_fd_pr__nfet_01v8__voff_diff_4 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_40 = {sky130_fd_pr__nfet_01v8__voff_diff_40 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_41 = {sky130_fd_pr__nfet_01v8__voff_diff_41 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_42 = {sky130_fd_pr__nfet_01v8__voff_diff_42 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_43 = {sky130_fd_pr__nfet_01v8__voff_diff_43 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_44 = {sky130_fd_pr__nfet_01v8__voff_diff_44 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_45 = {sky130_fd_pr__nfet_01v8__voff_diff_45 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_46 = {sky130_fd_pr__nfet_01v8__voff_diff_46 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_47 = {sky130_fd_pr__nfet_01v8__voff_diff_47 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_48 = {sky130_fd_pr__nfet_01v8__voff_diff_48 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_49 = {sky130_fd_pr__nfet_01v8__voff_diff_49 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_5 = {sky130_fd_pr__nfet_01v8__voff_diff_5 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_50 = {sky130_fd_pr__nfet_01v8__voff_diff_50 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_51 = {sky130_fd_pr__nfet_01v8__voff_diff_51 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_52 = {sky130_fd_pr__nfet_01v8__voff_diff_52 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_53 = {sky130_fd_pr__nfet_01v8__voff_diff_53 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_54 = {sky130_fd_pr__nfet_01v8__voff_diff_54 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_55 = {sky130_fd_pr__nfet_01v8__voff_diff_55 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_56 = {sky130_fd_pr__nfet_01v8__voff_diff_56 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_57 = {sky130_fd_pr__nfet_01v8__voff_diff_57 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_58 = {sky130_fd_pr__nfet_01v8__voff_diff_58 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_59 = {sky130_fd_pr__nfet_01v8__voff_diff_59 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_6 = {sky130_fd_pr__nfet_01v8__voff_diff_6 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_60 = {sky130_fd_pr__nfet_01v8__voff_diff_60 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_61 = {sky130_fd_pr__nfet_01v8__voff_diff_61 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_62 = {sky130_fd_pr__nfet_01v8__voff_diff_62 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_7 = {sky130_fd_pr__nfet_01v8__voff_diff_7 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_8 = {sky130_fd_pr__nfet_01v8__voff_diff_8 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__voff_diff_9 = {sky130_fd_pr__nfet_01v8__voff_diff_9 + k_nfet_voff_diff_cd*X_cd + k_nfet_voff_diff_damage*X_damage + k_nfet_voff_diff_eot*X_eot + k_nfet_voff_diff_act*X_act + k_nfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_0 = {sky130_fd_pr__nfet_01v8__vsat_diff_0 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_1 = {sky130_fd_pr__nfet_01v8__vsat_diff_1 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_10 = {sky130_fd_pr__nfet_01v8__vsat_diff_10 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_11 = {sky130_fd_pr__nfet_01v8__vsat_diff_11 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_12 = {sky130_fd_pr__nfet_01v8__vsat_diff_12 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_13 = {sky130_fd_pr__nfet_01v8__vsat_diff_13 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_14 = {sky130_fd_pr__nfet_01v8__vsat_diff_14 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_15 = {sky130_fd_pr__nfet_01v8__vsat_diff_15 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_16 = {sky130_fd_pr__nfet_01v8__vsat_diff_16 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_17 = {sky130_fd_pr__nfet_01v8__vsat_diff_17 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_18 = {sky130_fd_pr__nfet_01v8__vsat_diff_18 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_19 = {sky130_fd_pr__nfet_01v8__vsat_diff_19 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_2 = {sky130_fd_pr__nfet_01v8__vsat_diff_2 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_20 = {sky130_fd_pr__nfet_01v8__vsat_diff_20 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_21 = {sky130_fd_pr__nfet_01v8__vsat_diff_21 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_22 = {sky130_fd_pr__nfet_01v8__vsat_diff_22 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_23 = {sky130_fd_pr__nfet_01v8__vsat_diff_23 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_24 = {sky130_fd_pr__nfet_01v8__vsat_diff_24 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_25 = {sky130_fd_pr__nfet_01v8__vsat_diff_25 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_26 = {sky130_fd_pr__nfet_01v8__vsat_diff_26 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_27 = {sky130_fd_pr__nfet_01v8__vsat_diff_27 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_28 = {sky130_fd_pr__nfet_01v8__vsat_diff_28 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_29 = {sky130_fd_pr__nfet_01v8__vsat_diff_29 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_3 = {sky130_fd_pr__nfet_01v8__vsat_diff_3 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_30 = {sky130_fd_pr__nfet_01v8__vsat_diff_30 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_31 = {sky130_fd_pr__nfet_01v8__vsat_diff_31 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_32 = {sky130_fd_pr__nfet_01v8__vsat_diff_32 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_33 = {sky130_fd_pr__nfet_01v8__vsat_diff_33 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_34 = {sky130_fd_pr__nfet_01v8__vsat_diff_34 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_35 = {sky130_fd_pr__nfet_01v8__vsat_diff_35 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_36 = {sky130_fd_pr__nfet_01v8__vsat_diff_36 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_37 = {sky130_fd_pr__nfet_01v8__vsat_diff_37 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_38 = {sky130_fd_pr__nfet_01v8__vsat_diff_38 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_39 = {sky130_fd_pr__nfet_01v8__vsat_diff_39 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_4 = {sky130_fd_pr__nfet_01v8__vsat_diff_4 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_40 = {sky130_fd_pr__nfet_01v8__vsat_diff_40 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_41 = {sky130_fd_pr__nfet_01v8__vsat_diff_41 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_42 = {sky130_fd_pr__nfet_01v8__vsat_diff_42 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_43 = {sky130_fd_pr__nfet_01v8__vsat_diff_43 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_44 = {sky130_fd_pr__nfet_01v8__vsat_diff_44 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_45 = {sky130_fd_pr__nfet_01v8__vsat_diff_45 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_46 = {sky130_fd_pr__nfet_01v8__vsat_diff_46 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_47 = {sky130_fd_pr__nfet_01v8__vsat_diff_47 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_48 = {sky130_fd_pr__nfet_01v8__vsat_diff_48 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_49 = {sky130_fd_pr__nfet_01v8__vsat_diff_49 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_5 = {sky130_fd_pr__nfet_01v8__vsat_diff_5 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_50 = {sky130_fd_pr__nfet_01v8__vsat_diff_50 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_51 = {sky130_fd_pr__nfet_01v8__vsat_diff_51 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_52 = {sky130_fd_pr__nfet_01v8__vsat_diff_52 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_53 = {sky130_fd_pr__nfet_01v8__vsat_diff_53 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_54 = {sky130_fd_pr__nfet_01v8__vsat_diff_54 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_55 = {sky130_fd_pr__nfet_01v8__vsat_diff_55 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_56 = {sky130_fd_pr__nfet_01v8__vsat_diff_56 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_57 = {sky130_fd_pr__nfet_01v8__vsat_diff_57 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_58 = {sky130_fd_pr__nfet_01v8__vsat_diff_58 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_59 = {sky130_fd_pr__nfet_01v8__vsat_diff_59 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_6 = {sky130_fd_pr__nfet_01v8__vsat_diff_6 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_60 = {sky130_fd_pr__nfet_01v8__vsat_diff_60 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_61 = {sky130_fd_pr__nfet_01v8__vsat_diff_61 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_62 = {sky130_fd_pr__nfet_01v8__vsat_diff_62 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_7 = {sky130_fd_pr__nfet_01v8__vsat_diff_7 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_8 = {sky130_fd_pr__nfet_01v8__vsat_diff_8 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vsat_diff_9 = {sky130_fd_pr__nfet_01v8__vsat_diff_9 + k_nfet_vsat_diff_cd*X_cd + k_nfet_vsat_diff_damage*X_damage + k_nfet_vsat_diff_eot*X_eot + k_nfet_vsat_diff_act*X_act + k_nfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_0 = {sky130_fd_pr__nfet_01v8__vth0_diff_0 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_1 = {sky130_fd_pr__nfet_01v8__vth0_diff_1 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_10 = {sky130_fd_pr__nfet_01v8__vth0_diff_10 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_11 = {sky130_fd_pr__nfet_01v8__vth0_diff_11 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_12 = {sky130_fd_pr__nfet_01v8__vth0_diff_12 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_13 = {sky130_fd_pr__nfet_01v8__vth0_diff_13 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_14 = {sky130_fd_pr__nfet_01v8__vth0_diff_14 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_15 = {sky130_fd_pr__nfet_01v8__vth0_diff_15 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_16 = {sky130_fd_pr__nfet_01v8__vth0_diff_16 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_17 = {sky130_fd_pr__nfet_01v8__vth0_diff_17 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_18 = {sky130_fd_pr__nfet_01v8__vth0_diff_18 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_19 = {sky130_fd_pr__nfet_01v8__vth0_diff_19 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_2 = {sky130_fd_pr__nfet_01v8__vth0_diff_2 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_20 = {sky130_fd_pr__nfet_01v8__vth0_diff_20 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_21 = {sky130_fd_pr__nfet_01v8__vth0_diff_21 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_22 = {sky130_fd_pr__nfet_01v8__vth0_diff_22 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_23 = {sky130_fd_pr__nfet_01v8__vth0_diff_23 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_24 = {sky130_fd_pr__nfet_01v8__vth0_diff_24 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_25 = {sky130_fd_pr__nfet_01v8__vth0_diff_25 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_26 = {sky130_fd_pr__nfet_01v8__vth0_diff_26 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_27 = {sky130_fd_pr__nfet_01v8__vth0_diff_27 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_28 = {sky130_fd_pr__nfet_01v8__vth0_diff_28 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_29 = {sky130_fd_pr__nfet_01v8__vth0_diff_29 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_3 = {sky130_fd_pr__nfet_01v8__vth0_diff_3 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_30 = {sky130_fd_pr__nfet_01v8__vth0_diff_30 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_31 = {sky130_fd_pr__nfet_01v8__vth0_diff_31 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_32 = {sky130_fd_pr__nfet_01v8__vth0_diff_32 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_33 = {sky130_fd_pr__nfet_01v8__vth0_diff_33 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_34 = {sky130_fd_pr__nfet_01v8__vth0_diff_34 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_35 = {sky130_fd_pr__nfet_01v8__vth0_diff_35 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_36 = {sky130_fd_pr__nfet_01v8__vth0_diff_36 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_37 = {sky130_fd_pr__nfet_01v8__vth0_diff_37 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_38 = {sky130_fd_pr__nfet_01v8__vth0_diff_38 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_39 = {sky130_fd_pr__nfet_01v8__vth0_diff_39 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_4 = {sky130_fd_pr__nfet_01v8__vth0_diff_4 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_40 = {sky130_fd_pr__nfet_01v8__vth0_diff_40 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_41 = {sky130_fd_pr__nfet_01v8__vth0_diff_41 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_42 = {sky130_fd_pr__nfet_01v8__vth0_diff_42 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_43 = {sky130_fd_pr__nfet_01v8__vth0_diff_43 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_44 = {sky130_fd_pr__nfet_01v8__vth0_diff_44 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_45 = {sky130_fd_pr__nfet_01v8__vth0_diff_45 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_46 = {sky130_fd_pr__nfet_01v8__vth0_diff_46 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_47 = {sky130_fd_pr__nfet_01v8__vth0_diff_47 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_48 = {sky130_fd_pr__nfet_01v8__vth0_diff_48 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_49 = {sky130_fd_pr__nfet_01v8__vth0_diff_49 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_5 = {sky130_fd_pr__nfet_01v8__vth0_diff_5 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_50 = {sky130_fd_pr__nfet_01v8__vth0_diff_50 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_51 = {sky130_fd_pr__nfet_01v8__vth0_diff_51 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_52 = {sky130_fd_pr__nfet_01v8__vth0_diff_52 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_53 = {sky130_fd_pr__nfet_01v8__vth0_diff_53 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_54 = {sky130_fd_pr__nfet_01v8__vth0_diff_54 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_55 = {sky130_fd_pr__nfet_01v8__vth0_diff_55 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_56 = {sky130_fd_pr__nfet_01v8__vth0_diff_56 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_57 = {sky130_fd_pr__nfet_01v8__vth0_diff_57 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_58 = {sky130_fd_pr__nfet_01v8__vth0_diff_58 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_59 = {sky130_fd_pr__nfet_01v8__vth0_diff_59 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_6 = {sky130_fd_pr__nfet_01v8__vth0_diff_6 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_60 = {sky130_fd_pr__nfet_01v8__vth0_diff_60 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_61 = {sky130_fd_pr__nfet_01v8__vth0_diff_61 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_62 = {sky130_fd_pr__nfet_01v8__vth0_diff_62 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_7 = {sky130_fd_pr__nfet_01v8__vth0_diff_7 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_8 = {sky130_fd_pr__nfet_01v8__vth0_diff_8 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__nfet_01v8__vth0_diff_9 = {sky130_fd_pr__nfet_01v8__vth0_diff_9 + k_nfet_vth0_diff_cd*X_cd + k_nfet_vth0_diff_damage*X_damage + k_nfet_vth0_diff_eot*X_eot + k_nfet_vth0_diff_act*X_act + k_nfet_vth0_diff_rc*X_rc}

* PFET equations
.param sky130_fd_pr__pfet_01v8__ajunction_mult = {sky130_fd_pr__pfet_01v8__ajunction_mult*(1 + k_pfet_ajunction_mult_cd*X_cd + k_pfet_ajunction_mult_damage*X_damage + k_pfet_ajunction_mult_eot*X_eot + k_pfet_ajunction_mult_act*X_act + k_pfet_ajunction_mult_rc*X_rc)}
.param sky130_fd_pr__pfet_01v8__dlc_diff = {sky130_fd_pr__pfet_01v8__dlc_diff + k_pfet_dlc_diff_cd*X_cd + k_pfet_dlc_diff_damage*X_damage + k_pfet_dlc_diff_eot*X_eot + k_pfet_dlc_diff_act*X_act + k_pfet_dlc_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__dwc_diff = {sky130_fd_pr__pfet_01v8__dwc_diff + k_pfet_dwc_diff_cd*X_cd + k_pfet_dwc_diff_damage*X_damage + k_pfet_dwc_diff_eot*X_eot + k_pfet_dwc_diff_act*X_act + k_pfet_dwc_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__lint_diff = {sky130_fd_pr__pfet_01v8__lint_diff + k_pfet_lint_diff_cd*X_cd + k_pfet_lint_diff_damage*X_damage + k_pfet_lint_diff_eot*X_eot + k_pfet_lint_diff_act*X_act + k_pfet_lint_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__overlap_mult = {sky130_fd_pr__pfet_01v8__overlap_mult*(1 + k_pfet_overlap_mult_cd*X_cd + k_pfet_overlap_mult_damage*X_damage + k_pfet_overlap_mult_eot*X_eot + k_pfet_overlap_mult_act*X_act + k_pfet_overlap_mult_rc*X_rc)}
.param sky130_fd_pr__pfet_01v8__pjunction_mult = {sky130_fd_pr__pfet_01v8__pjunction_mult*(1 + k_pfet_pjunction_mult_cd*X_cd + k_pfet_pjunction_mult_damage*X_damage + k_pfet_pjunction_mult_eot*X_eot + k_pfet_pjunction_mult_act*X_act + k_pfet_pjunction_mult_rc*X_rc)}
.param sky130_fd_pr__pfet_01v8__rshp_mult = {sky130_fd_pr__pfet_01v8__rshp_mult*(1 + k_pfet_rshp_mult_cd*X_cd + k_pfet_rshp_mult_damage*X_damage + k_pfet_rshp_mult_eot*X_eot + k_pfet_rshp_mult_act*X_act + k_pfet_rshp_mult_rc*X_rc)}
.param sky130_fd_pr__pfet_01v8__toxe_mult = {sky130_fd_pr__pfet_01v8__toxe_mult*(1 + k_pfet_toxe_mult_cd*X_cd + k_pfet_toxe_mult_damage*X_damage + k_pfet_toxe_mult_eot*X_eot + k_pfet_toxe_mult_act*X_act + k_pfet_toxe_mult_rc*X_rc)}
.param sky130_fd_pr__pfet_01v8__wint_diff = {sky130_fd_pr__pfet_01v8__wint_diff + k_pfet_wint_diff_cd*X_cd + k_pfet_wint_diff_damage*X_damage + k_pfet_wint_diff_eot*X_eot + k_pfet_wint_diff_act*X_act + k_pfet_wint_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_0 = {sky130_fd_pr__pfet_01v8__a0_diff_0 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_1 = {sky130_fd_pr__pfet_01v8__a0_diff_1 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_10 = {sky130_fd_pr__pfet_01v8__a0_diff_10 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_11 = {sky130_fd_pr__pfet_01v8__a0_diff_11 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_12 = {sky130_fd_pr__pfet_01v8__a0_diff_12 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_13 = {sky130_fd_pr__pfet_01v8__a0_diff_13 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_14 = {sky130_fd_pr__pfet_01v8__a0_diff_14 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_15 = {sky130_fd_pr__pfet_01v8__a0_diff_15 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_16 = {sky130_fd_pr__pfet_01v8__a0_diff_16 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_17 = {sky130_fd_pr__pfet_01v8__a0_diff_17 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_18 = {sky130_fd_pr__pfet_01v8__a0_diff_18 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_19 = {sky130_fd_pr__pfet_01v8__a0_diff_19 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_2 = {sky130_fd_pr__pfet_01v8__a0_diff_2 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_20 = {sky130_fd_pr__pfet_01v8__a0_diff_20 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_21 = {sky130_fd_pr__pfet_01v8__a0_diff_21 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_22 = {sky130_fd_pr__pfet_01v8__a0_diff_22 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_23 = {sky130_fd_pr__pfet_01v8__a0_diff_23 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_24 = {sky130_fd_pr__pfet_01v8__a0_diff_24 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_25 = {sky130_fd_pr__pfet_01v8__a0_diff_25 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_26 = {sky130_fd_pr__pfet_01v8__a0_diff_26 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_27 = {sky130_fd_pr__pfet_01v8__a0_diff_27 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_28 = {sky130_fd_pr__pfet_01v8__a0_diff_28 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_29 = {sky130_fd_pr__pfet_01v8__a0_diff_29 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_3 = {sky130_fd_pr__pfet_01v8__a0_diff_3 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_30 = {sky130_fd_pr__pfet_01v8__a0_diff_30 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_31 = {sky130_fd_pr__pfet_01v8__a0_diff_31 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_32 = {sky130_fd_pr__pfet_01v8__a0_diff_32 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_33 = {sky130_fd_pr__pfet_01v8__a0_diff_33 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_34 = {sky130_fd_pr__pfet_01v8__a0_diff_34 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_35 = {sky130_fd_pr__pfet_01v8__a0_diff_35 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_36 = {sky130_fd_pr__pfet_01v8__a0_diff_36 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_37 = {sky130_fd_pr__pfet_01v8__a0_diff_37 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_38 = {sky130_fd_pr__pfet_01v8__a0_diff_38 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_39 = {sky130_fd_pr__pfet_01v8__a0_diff_39 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_4 = {sky130_fd_pr__pfet_01v8__a0_diff_4 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_40 = {sky130_fd_pr__pfet_01v8__a0_diff_40 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_41 = {sky130_fd_pr__pfet_01v8__a0_diff_41 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_42 = {sky130_fd_pr__pfet_01v8__a0_diff_42 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_43 = {sky130_fd_pr__pfet_01v8__a0_diff_43 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_44 = {sky130_fd_pr__pfet_01v8__a0_diff_44 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_45 = {sky130_fd_pr__pfet_01v8__a0_diff_45 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_46 = {sky130_fd_pr__pfet_01v8__a0_diff_46 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_47 = {sky130_fd_pr__pfet_01v8__a0_diff_47 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_48 = {sky130_fd_pr__pfet_01v8__a0_diff_48 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_49 = {sky130_fd_pr__pfet_01v8__a0_diff_49 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_5 = {sky130_fd_pr__pfet_01v8__a0_diff_5 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_50 = {sky130_fd_pr__pfet_01v8__a0_diff_50 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_51 = {sky130_fd_pr__pfet_01v8__a0_diff_51 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_6 = {sky130_fd_pr__pfet_01v8__a0_diff_6 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_7 = {sky130_fd_pr__pfet_01v8__a0_diff_7 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_8 = {sky130_fd_pr__pfet_01v8__a0_diff_8 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__a0_diff_9 = {sky130_fd_pr__pfet_01v8__a0_diff_9 + k_pfet_a0_diff_cd*X_cd + k_pfet_a0_diff_damage*X_damage + k_pfet_a0_diff_eot*X_eot + k_pfet_a0_diff_act*X_act + k_pfet_a0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_0 = {sky130_fd_pr__pfet_01v8__agidl_diff_0 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_1 = {sky130_fd_pr__pfet_01v8__agidl_diff_1 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_10 = {sky130_fd_pr__pfet_01v8__agidl_diff_10 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_11 = {sky130_fd_pr__pfet_01v8__agidl_diff_11 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_12 = {sky130_fd_pr__pfet_01v8__agidl_diff_12 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_13 = {sky130_fd_pr__pfet_01v8__agidl_diff_13 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_14 = {sky130_fd_pr__pfet_01v8__agidl_diff_14 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_15 = {sky130_fd_pr__pfet_01v8__agidl_diff_15 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_16 = {sky130_fd_pr__pfet_01v8__agidl_diff_16 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_17 = {sky130_fd_pr__pfet_01v8__agidl_diff_17 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_18 = {sky130_fd_pr__pfet_01v8__agidl_diff_18 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_19 = {sky130_fd_pr__pfet_01v8__agidl_diff_19 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_2 = {sky130_fd_pr__pfet_01v8__agidl_diff_2 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_20 = {sky130_fd_pr__pfet_01v8__agidl_diff_20 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_21 = {sky130_fd_pr__pfet_01v8__agidl_diff_21 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_22 = {sky130_fd_pr__pfet_01v8__agidl_diff_22 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_23 = {sky130_fd_pr__pfet_01v8__agidl_diff_23 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_24 = {sky130_fd_pr__pfet_01v8__agidl_diff_24 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_25 = {sky130_fd_pr__pfet_01v8__agidl_diff_25 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_26 = {sky130_fd_pr__pfet_01v8__agidl_diff_26 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_27 = {sky130_fd_pr__pfet_01v8__agidl_diff_27 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_28 = {sky130_fd_pr__pfet_01v8__agidl_diff_28 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_29 = {sky130_fd_pr__pfet_01v8__agidl_diff_29 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_3 = {sky130_fd_pr__pfet_01v8__agidl_diff_3 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_30 = {sky130_fd_pr__pfet_01v8__agidl_diff_30 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_31 = {sky130_fd_pr__pfet_01v8__agidl_diff_31 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_32 = {sky130_fd_pr__pfet_01v8__agidl_diff_32 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_33 = {sky130_fd_pr__pfet_01v8__agidl_diff_33 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_34 = {sky130_fd_pr__pfet_01v8__agidl_diff_34 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_35 = {sky130_fd_pr__pfet_01v8__agidl_diff_35 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_36 = {sky130_fd_pr__pfet_01v8__agidl_diff_36 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_37 = {sky130_fd_pr__pfet_01v8__agidl_diff_37 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_38 = {sky130_fd_pr__pfet_01v8__agidl_diff_38 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_39 = {sky130_fd_pr__pfet_01v8__agidl_diff_39 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_4 = {sky130_fd_pr__pfet_01v8__agidl_diff_4 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_40 = {sky130_fd_pr__pfet_01v8__agidl_diff_40 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_41 = {sky130_fd_pr__pfet_01v8__agidl_diff_41 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_42 = {sky130_fd_pr__pfet_01v8__agidl_diff_42 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_43 = {sky130_fd_pr__pfet_01v8__agidl_diff_43 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_44 = {sky130_fd_pr__pfet_01v8__agidl_diff_44 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_45 = {sky130_fd_pr__pfet_01v8__agidl_diff_45 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_46 = {sky130_fd_pr__pfet_01v8__agidl_diff_46 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_47 = {sky130_fd_pr__pfet_01v8__agidl_diff_47 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_48 = {sky130_fd_pr__pfet_01v8__agidl_diff_48 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_49 = {sky130_fd_pr__pfet_01v8__agidl_diff_49 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_5 = {sky130_fd_pr__pfet_01v8__agidl_diff_5 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_50 = {sky130_fd_pr__pfet_01v8__agidl_diff_50 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_51 = {sky130_fd_pr__pfet_01v8__agidl_diff_51 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_6 = {sky130_fd_pr__pfet_01v8__agidl_diff_6 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_7 = {sky130_fd_pr__pfet_01v8__agidl_diff_7 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_8 = {sky130_fd_pr__pfet_01v8__agidl_diff_8 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__agidl_diff_9 = {sky130_fd_pr__pfet_01v8__agidl_diff_9 + k_pfet_agidl_diff_cd*X_cd + k_pfet_agidl_diff_damage*X_damage + k_pfet_agidl_diff_eot*X_eot + k_pfet_agidl_diff_act*X_act + k_pfet_agidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_0 = {sky130_fd_pr__pfet_01v8__ags_diff_0 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_1 = {sky130_fd_pr__pfet_01v8__ags_diff_1 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_10 = {sky130_fd_pr__pfet_01v8__ags_diff_10 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_11 = {sky130_fd_pr__pfet_01v8__ags_diff_11 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_12 = {sky130_fd_pr__pfet_01v8__ags_diff_12 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_13 = {sky130_fd_pr__pfet_01v8__ags_diff_13 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_14 = {sky130_fd_pr__pfet_01v8__ags_diff_14 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_15 = {sky130_fd_pr__pfet_01v8__ags_diff_15 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_16 = {sky130_fd_pr__pfet_01v8__ags_diff_16 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_17 = {sky130_fd_pr__pfet_01v8__ags_diff_17 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_18 = {sky130_fd_pr__pfet_01v8__ags_diff_18 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_19 = {sky130_fd_pr__pfet_01v8__ags_diff_19 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_2 = {sky130_fd_pr__pfet_01v8__ags_diff_2 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_20 = {sky130_fd_pr__pfet_01v8__ags_diff_20 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_21 = {sky130_fd_pr__pfet_01v8__ags_diff_21 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_22 = {sky130_fd_pr__pfet_01v8__ags_diff_22 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_23 = {sky130_fd_pr__pfet_01v8__ags_diff_23 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_24 = {sky130_fd_pr__pfet_01v8__ags_diff_24 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_25 = {sky130_fd_pr__pfet_01v8__ags_diff_25 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_26 = {sky130_fd_pr__pfet_01v8__ags_diff_26 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_27 = {sky130_fd_pr__pfet_01v8__ags_diff_27 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_28 = {sky130_fd_pr__pfet_01v8__ags_diff_28 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_29 = {sky130_fd_pr__pfet_01v8__ags_diff_29 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_3 = {sky130_fd_pr__pfet_01v8__ags_diff_3 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_30 = {sky130_fd_pr__pfet_01v8__ags_diff_30 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_31 = {sky130_fd_pr__pfet_01v8__ags_diff_31 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_32 = {sky130_fd_pr__pfet_01v8__ags_diff_32 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_33 = {sky130_fd_pr__pfet_01v8__ags_diff_33 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_34 = {sky130_fd_pr__pfet_01v8__ags_diff_34 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_35 = {sky130_fd_pr__pfet_01v8__ags_diff_35 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_36 = {sky130_fd_pr__pfet_01v8__ags_diff_36 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_37 = {sky130_fd_pr__pfet_01v8__ags_diff_37 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_38 = {sky130_fd_pr__pfet_01v8__ags_diff_38 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_39 = {sky130_fd_pr__pfet_01v8__ags_diff_39 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_4 = {sky130_fd_pr__pfet_01v8__ags_diff_4 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_40 = {sky130_fd_pr__pfet_01v8__ags_diff_40 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_41 = {sky130_fd_pr__pfet_01v8__ags_diff_41 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_42 = {sky130_fd_pr__pfet_01v8__ags_diff_42 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_43 = {sky130_fd_pr__pfet_01v8__ags_diff_43 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_44 = {sky130_fd_pr__pfet_01v8__ags_diff_44 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_45 = {sky130_fd_pr__pfet_01v8__ags_diff_45 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_46 = {sky130_fd_pr__pfet_01v8__ags_diff_46 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_47 = {sky130_fd_pr__pfet_01v8__ags_diff_47 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_48 = {sky130_fd_pr__pfet_01v8__ags_diff_48 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_49 = {sky130_fd_pr__pfet_01v8__ags_diff_49 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_5 = {sky130_fd_pr__pfet_01v8__ags_diff_5 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_50 = {sky130_fd_pr__pfet_01v8__ags_diff_50 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_51 = {sky130_fd_pr__pfet_01v8__ags_diff_51 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_6 = {sky130_fd_pr__pfet_01v8__ags_diff_6 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_7 = {sky130_fd_pr__pfet_01v8__ags_diff_7 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_8 = {sky130_fd_pr__pfet_01v8__ags_diff_8 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ags_diff_9 = {sky130_fd_pr__pfet_01v8__ags_diff_9 + k_pfet_ags_diff_cd*X_cd + k_pfet_ags_diff_damage*X_damage + k_pfet_ags_diff_eot*X_eot + k_pfet_ags_diff_act*X_act + k_pfet_ags_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_0 = {sky130_fd_pr__pfet_01v8__b0_diff_0 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_1 = {sky130_fd_pr__pfet_01v8__b0_diff_1 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_10 = {sky130_fd_pr__pfet_01v8__b0_diff_10 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_11 = {sky130_fd_pr__pfet_01v8__b0_diff_11 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_12 = {sky130_fd_pr__pfet_01v8__b0_diff_12 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_13 = {sky130_fd_pr__pfet_01v8__b0_diff_13 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_14 = {sky130_fd_pr__pfet_01v8__b0_diff_14 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_15 = {sky130_fd_pr__pfet_01v8__b0_diff_15 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_16 = {sky130_fd_pr__pfet_01v8__b0_diff_16 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_17 = {sky130_fd_pr__pfet_01v8__b0_diff_17 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_18 = {sky130_fd_pr__pfet_01v8__b0_diff_18 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_19 = {sky130_fd_pr__pfet_01v8__b0_diff_19 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_2 = {sky130_fd_pr__pfet_01v8__b0_diff_2 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_20 = {sky130_fd_pr__pfet_01v8__b0_diff_20 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_21 = {sky130_fd_pr__pfet_01v8__b0_diff_21 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_22 = {sky130_fd_pr__pfet_01v8__b0_diff_22 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_23 = {sky130_fd_pr__pfet_01v8__b0_diff_23 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_24 = {sky130_fd_pr__pfet_01v8__b0_diff_24 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_25 = {sky130_fd_pr__pfet_01v8__b0_diff_25 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_26 = {sky130_fd_pr__pfet_01v8__b0_diff_26 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_27 = {sky130_fd_pr__pfet_01v8__b0_diff_27 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_28 = {sky130_fd_pr__pfet_01v8__b0_diff_28 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_29 = {sky130_fd_pr__pfet_01v8__b0_diff_29 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_3 = {sky130_fd_pr__pfet_01v8__b0_diff_3 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_30 = {sky130_fd_pr__pfet_01v8__b0_diff_30 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_31 = {sky130_fd_pr__pfet_01v8__b0_diff_31 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_32 = {sky130_fd_pr__pfet_01v8__b0_diff_32 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_33 = {sky130_fd_pr__pfet_01v8__b0_diff_33 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_34 = {sky130_fd_pr__pfet_01v8__b0_diff_34 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_35 = {sky130_fd_pr__pfet_01v8__b0_diff_35 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_36 = {sky130_fd_pr__pfet_01v8__b0_diff_36 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_37 = {sky130_fd_pr__pfet_01v8__b0_diff_37 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_38 = {sky130_fd_pr__pfet_01v8__b0_diff_38 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_39 = {sky130_fd_pr__pfet_01v8__b0_diff_39 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_4 = {sky130_fd_pr__pfet_01v8__b0_diff_4 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_40 = {sky130_fd_pr__pfet_01v8__b0_diff_40 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_41 = {sky130_fd_pr__pfet_01v8__b0_diff_41 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_42 = {sky130_fd_pr__pfet_01v8__b0_diff_42 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_43 = {sky130_fd_pr__pfet_01v8__b0_diff_43 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_44 = {sky130_fd_pr__pfet_01v8__b0_diff_44 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_45 = {sky130_fd_pr__pfet_01v8__b0_diff_45 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_46 = {sky130_fd_pr__pfet_01v8__b0_diff_46 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_47 = {sky130_fd_pr__pfet_01v8__b0_diff_47 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_48 = {sky130_fd_pr__pfet_01v8__b0_diff_48 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_49 = {sky130_fd_pr__pfet_01v8__b0_diff_49 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_5 = {sky130_fd_pr__pfet_01v8__b0_diff_5 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_50 = {sky130_fd_pr__pfet_01v8__b0_diff_50 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_51 = {sky130_fd_pr__pfet_01v8__b0_diff_51 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_6 = {sky130_fd_pr__pfet_01v8__b0_diff_6 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_7 = {sky130_fd_pr__pfet_01v8__b0_diff_7 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_8 = {sky130_fd_pr__pfet_01v8__b0_diff_8 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b0_diff_9 = {sky130_fd_pr__pfet_01v8__b0_diff_9 + k_pfet_b0_diff_cd*X_cd + k_pfet_b0_diff_damage*X_damage + k_pfet_b0_diff_eot*X_eot + k_pfet_b0_diff_act*X_act + k_pfet_b0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_0 = {sky130_fd_pr__pfet_01v8__b1_diff_0 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_1 = {sky130_fd_pr__pfet_01v8__b1_diff_1 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_10 = {sky130_fd_pr__pfet_01v8__b1_diff_10 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_11 = {sky130_fd_pr__pfet_01v8__b1_diff_11 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_12 = {sky130_fd_pr__pfet_01v8__b1_diff_12 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_13 = {sky130_fd_pr__pfet_01v8__b1_diff_13 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_14 = {sky130_fd_pr__pfet_01v8__b1_diff_14 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_15 = {sky130_fd_pr__pfet_01v8__b1_diff_15 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_16 = {sky130_fd_pr__pfet_01v8__b1_diff_16 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_17 = {sky130_fd_pr__pfet_01v8__b1_diff_17 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_18 = {sky130_fd_pr__pfet_01v8__b1_diff_18 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_19 = {sky130_fd_pr__pfet_01v8__b1_diff_19 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_2 = {sky130_fd_pr__pfet_01v8__b1_diff_2 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_20 = {sky130_fd_pr__pfet_01v8__b1_diff_20 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_21 = {sky130_fd_pr__pfet_01v8__b1_diff_21 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_22 = {sky130_fd_pr__pfet_01v8__b1_diff_22 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_23 = {sky130_fd_pr__pfet_01v8__b1_diff_23 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_24 = {sky130_fd_pr__pfet_01v8__b1_diff_24 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_25 = {sky130_fd_pr__pfet_01v8__b1_diff_25 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_26 = {sky130_fd_pr__pfet_01v8__b1_diff_26 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_27 = {sky130_fd_pr__pfet_01v8__b1_diff_27 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_28 = {sky130_fd_pr__pfet_01v8__b1_diff_28 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_29 = {sky130_fd_pr__pfet_01v8__b1_diff_29 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_3 = {sky130_fd_pr__pfet_01v8__b1_diff_3 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_30 = {sky130_fd_pr__pfet_01v8__b1_diff_30 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_31 = {sky130_fd_pr__pfet_01v8__b1_diff_31 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_32 = {sky130_fd_pr__pfet_01v8__b1_diff_32 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_33 = {sky130_fd_pr__pfet_01v8__b1_diff_33 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_34 = {sky130_fd_pr__pfet_01v8__b1_diff_34 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_35 = {sky130_fd_pr__pfet_01v8__b1_diff_35 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_36 = {sky130_fd_pr__pfet_01v8__b1_diff_36 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_37 = {sky130_fd_pr__pfet_01v8__b1_diff_37 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_38 = {sky130_fd_pr__pfet_01v8__b1_diff_38 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_39 = {sky130_fd_pr__pfet_01v8__b1_diff_39 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_4 = {sky130_fd_pr__pfet_01v8__b1_diff_4 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_40 = {sky130_fd_pr__pfet_01v8__b1_diff_40 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_41 = {sky130_fd_pr__pfet_01v8__b1_diff_41 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_42 = {sky130_fd_pr__pfet_01v8__b1_diff_42 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_43 = {sky130_fd_pr__pfet_01v8__b1_diff_43 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_44 = {sky130_fd_pr__pfet_01v8__b1_diff_44 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_45 = {sky130_fd_pr__pfet_01v8__b1_diff_45 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_46 = {sky130_fd_pr__pfet_01v8__b1_diff_46 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_47 = {sky130_fd_pr__pfet_01v8__b1_diff_47 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_48 = {sky130_fd_pr__pfet_01v8__b1_diff_48 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_49 = {sky130_fd_pr__pfet_01v8__b1_diff_49 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_5 = {sky130_fd_pr__pfet_01v8__b1_diff_5 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_50 = {sky130_fd_pr__pfet_01v8__b1_diff_50 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_51 = {sky130_fd_pr__pfet_01v8__b1_diff_51 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_6 = {sky130_fd_pr__pfet_01v8__b1_diff_6 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_7 = {sky130_fd_pr__pfet_01v8__b1_diff_7 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_8 = {sky130_fd_pr__pfet_01v8__b1_diff_8 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__b1_diff_9 = {sky130_fd_pr__pfet_01v8__b1_diff_9 + k_pfet_b1_diff_cd*X_cd + k_pfet_b1_diff_damage*X_damage + k_pfet_b1_diff_eot*X_eot + k_pfet_b1_diff_act*X_act + k_pfet_b1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_0 = {sky130_fd_pr__pfet_01v8__bgidl_diff_0 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_1 = {sky130_fd_pr__pfet_01v8__bgidl_diff_1 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_10 = {sky130_fd_pr__pfet_01v8__bgidl_diff_10 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_11 = {sky130_fd_pr__pfet_01v8__bgidl_diff_11 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_12 = {sky130_fd_pr__pfet_01v8__bgidl_diff_12 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_13 = {sky130_fd_pr__pfet_01v8__bgidl_diff_13 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_14 = {sky130_fd_pr__pfet_01v8__bgidl_diff_14 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_15 = {sky130_fd_pr__pfet_01v8__bgidl_diff_15 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_16 = {sky130_fd_pr__pfet_01v8__bgidl_diff_16 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_17 = {sky130_fd_pr__pfet_01v8__bgidl_diff_17 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_18 = {sky130_fd_pr__pfet_01v8__bgidl_diff_18 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_19 = {sky130_fd_pr__pfet_01v8__bgidl_diff_19 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_2 = {sky130_fd_pr__pfet_01v8__bgidl_diff_2 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_20 = {sky130_fd_pr__pfet_01v8__bgidl_diff_20 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_21 = {sky130_fd_pr__pfet_01v8__bgidl_diff_21 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_22 = {sky130_fd_pr__pfet_01v8__bgidl_diff_22 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_23 = {sky130_fd_pr__pfet_01v8__bgidl_diff_23 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_24 = {sky130_fd_pr__pfet_01v8__bgidl_diff_24 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_25 = {sky130_fd_pr__pfet_01v8__bgidl_diff_25 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_26 = {sky130_fd_pr__pfet_01v8__bgidl_diff_26 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_27 = {sky130_fd_pr__pfet_01v8__bgidl_diff_27 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_28 = {sky130_fd_pr__pfet_01v8__bgidl_diff_28 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_29 = {sky130_fd_pr__pfet_01v8__bgidl_diff_29 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_3 = {sky130_fd_pr__pfet_01v8__bgidl_diff_3 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_30 = {sky130_fd_pr__pfet_01v8__bgidl_diff_30 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_31 = {sky130_fd_pr__pfet_01v8__bgidl_diff_31 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_32 = {sky130_fd_pr__pfet_01v8__bgidl_diff_32 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_33 = {sky130_fd_pr__pfet_01v8__bgidl_diff_33 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_34 = {sky130_fd_pr__pfet_01v8__bgidl_diff_34 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_35 = {sky130_fd_pr__pfet_01v8__bgidl_diff_35 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_36 = {sky130_fd_pr__pfet_01v8__bgidl_diff_36 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_37 = {sky130_fd_pr__pfet_01v8__bgidl_diff_37 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_38 = {sky130_fd_pr__pfet_01v8__bgidl_diff_38 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_39 = {sky130_fd_pr__pfet_01v8__bgidl_diff_39 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_4 = {sky130_fd_pr__pfet_01v8__bgidl_diff_4 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_40 = {sky130_fd_pr__pfet_01v8__bgidl_diff_40 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_41 = {sky130_fd_pr__pfet_01v8__bgidl_diff_41 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_42 = {sky130_fd_pr__pfet_01v8__bgidl_diff_42 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_43 = {sky130_fd_pr__pfet_01v8__bgidl_diff_43 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_44 = {sky130_fd_pr__pfet_01v8__bgidl_diff_44 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_45 = {sky130_fd_pr__pfet_01v8__bgidl_diff_45 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_46 = {sky130_fd_pr__pfet_01v8__bgidl_diff_46 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_47 = {sky130_fd_pr__pfet_01v8__bgidl_diff_47 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_48 = {sky130_fd_pr__pfet_01v8__bgidl_diff_48 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_49 = {sky130_fd_pr__pfet_01v8__bgidl_diff_49 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_5 = {sky130_fd_pr__pfet_01v8__bgidl_diff_5 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_50 = {sky130_fd_pr__pfet_01v8__bgidl_diff_50 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_51 = {sky130_fd_pr__pfet_01v8__bgidl_diff_51 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_6 = {sky130_fd_pr__pfet_01v8__bgidl_diff_6 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_7 = {sky130_fd_pr__pfet_01v8__bgidl_diff_7 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_8 = {sky130_fd_pr__pfet_01v8__bgidl_diff_8 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__bgidl_diff_9 = {sky130_fd_pr__pfet_01v8__bgidl_diff_9 + k_pfet_bgidl_diff_cd*X_cd + k_pfet_bgidl_diff_damage*X_damage + k_pfet_bgidl_diff_eot*X_eot + k_pfet_bgidl_diff_act*X_act + k_pfet_bgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_0 = {sky130_fd_pr__pfet_01v8__cgidl_diff_0 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_1 = {sky130_fd_pr__pfet_01v8__cgidl_diff_1 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_10 = {sky130_fd_pr__pfet_01v8__cgidl_diff_10 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_11 = {sky130_fd_pr__pfet_01v8__cgidl_diff_11 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_12 = {sky130_fd_pr__pfet_01v8__cgidl_diff_12 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_13 = {sky130_fd_pr__pfet_01v8__cgidl_diff_13 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_14 = {sky130_fd_pr__pfet_01v8__cgidl_diff_14 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_15 = {sky130_fd_pr__pfet_01v8__cgidl_diff_15 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_16 = {sky130_fd_pr__pfet_01v8__cgidl_diff_16 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_17 = {sky130_fd_pr__pfet_01v8__cgidl_diff_17 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_18 = {sky130_fd_pr__pfet_01v8__cgidl_diff_18 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_19 = {sky130_fd_pr__pfet_01v8__cgidl_diff_19 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_2 = {sky130_fd_pr__pfet_01v8__cgidl_diff_2 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_20 = {sky130_fd_pr__pfet_01v8__cgidl_diff_20 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_21 = {sky130_fd_pr__pfet_01v8__cgidl_diff_21 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_22 = {sky130_fd_pr__pfet_01v8__cgidl_diff_22 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_23 = {sky130_fd_pr__pfet_01v8__cgidl_diff_23 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_24 = {sky130_fd_pr__pfet_01v8__cgidl_diff_24 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_25 = {sky130_fd_pr__pfet_01v8__cgidl_diff_25 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_26 = {sky130_fd_pr__pfet_01v8__cgidl_diff_26 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_27 = {sky130_fd_pr__pfet_01v8__cgidl_diff_27 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_28 = {sky130_fd_pr__pfet_01v8__cgidl_diff_28 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_29 = {sky130_fd_pr__pfet_01v8__cgidl_diff_29 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_3 = {sky130_fd_pr__pfet_01v8__cgidl_diff_3 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_30 = {sky130_fd_pr__pfet_01v8__cgidl_diff_30 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_31 = {sky130_fd_pr__pfet_01v8__cgidl_diff_31 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_32 = {sky130_fd_pr__pfet_01v8__cgidl_diff_32 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_33 = {sky130_fd_pr__pfet_01v8__cgidl_diff_33 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_34 = {sky130_fd_pr__pfet_01v8__cgidl_diff_34 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_35 = {sky130_fd_pr__pfet_01v8__cgidl_diff_35 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_36 = {sky130_fd_pr__pfet_01v8__cgidl_diff_36 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_37 = {sky130_fd_pr__pfet_01v8__cgidl_diff_37 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_38 = {sky130_fd_pr__pfet_01v8__cgidl_diff_38 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_39 = {sky130_fd_pr__pfet_01v8__cgidl_diff_39 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_4 = {sky130_fd_pr__pfet_01v8__cgidl_diff_4 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_40 = {sky130_fd_pr__pfet_01v8__cgidl_diff_40 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_41 = {sky130_fd_pr__pfet_01v8__cgidl_diff_41 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_42 = {sky130_fd_pr__pfet_01v8__cgidl_diff_42 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_43 = {sky130_fd_pr__pfet_01v8__cgidl_diff_43 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_44 = {sky130_fd_pr__pfet_01v8__cgidl_diff_44 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_45 = {sky130_fd_pr__pfet_01v8__cgidl_diff_45 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_46 = {sky130_fd_pr__pfet_01v8__cgidl_diff_46 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_47 = {sky130_fd_pr__pfet_01v8__cgidl_diff_47 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_48 = {sky130_fd_pr__pfet_01v8__cgidl_diff_48 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_49 = {sky130_fd_pr__pfet_01v8__cgidl_diff_49 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_5 = {sky130_fd_pr__pfet_01v8__cgidl_diff_5 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_50 = {sky130_fd_pr__pfet_01v8__cgidl_diff_50 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_51 = {sky130_fd_pr__pfet_01v8__cgidl_diff_51 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_6 = {sky130_fd_pr__pfet_01v8__cgidl_diff_6 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_7 = {sky130_fd_pr__pfet_01v8__cgidl_diff_7 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_8 = {sky130_fd_pr__pfet_01v8__cgidl_diff_8 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__cgidl_diff_9 = {sky130_fd_pr__pfet_01v8__cgidl_diff_9 + k_pfet_cgidl_diff_cd*X_cd + k_pfet_cgidl_diff_damage*X_damage + k_pfet_cgidl_diff_eot*X_eot + k_pfet_cgidl_diff_act*X_act + k_pfet_cgidl_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_0 = {sky130_fd_pr__pfet_01v8__eta0_diff_0 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_1 = {sky130_fd_pr__pfet_01v8__eta0_diff_1 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_10 = {sky130_fd_pr__pfet_01v8__eta0_diff_10 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_11 = {sky130_fd_pr__pfet_01v8__eta0_diff_11 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_12 = {sky130_fd_pr__pfet_01v8__eta0_diff_12 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_13 = {sky130_fd_pr__pfet_01v8__eta0_diff_13 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_14 = {sky130_fd_pr__pfet_01v8__eta0_diff_14 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_15 = {sky130_fd_pr__pfet_01v8__eta0_diff_15 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_16 = {sky130_fd_pr__pfet_01v8__eta0_diff_16 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_17 = {sky130_fd_pr__pfet_01v8__eta0_diff_17 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_18 = {sky130_fd_pr__pfet_01v8__eta0_diff_18 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_19 = {sky130_fd_pr__pfet_01v8__eta0_diff_19 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_2 = {sky130_fd_pr__pfet_01v8__eta0_diff_2 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_20 = {sky130_fd_pr__pfet_01v8__eta0_diff_20 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_21 = {sky130_fd_pr__pfet_01v8__eta0_diff_21 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_22 = {sky130_fd_pr__pfet_01v8__eta0_diff_22 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_23 = {sky130_fd_pr__pfet_01v8__eta0_diff_23 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_24 = {sky130_fd_pr__pfet_01v8__eta0_diff_24 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_25 = {sky130_fd_pr__pfet_01v8__eta0_diff_25 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_26 = {sky130_fd_pr__pfet_01v8__eta0_diff_26 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_27 = {sky130_fd_pr__pfet_01v8__eta0_diff_27 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_28 = {sky130_fd_pr__pfet_01v8__eta0_diff_28 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_29 = {sky130_fd_pr__pfet_01v8__eta0_diff_29 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_3 = {sky130_fd_pr__pfet_01v8__eta0_diff_3 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_30 = {sky130_fd_pr__pfet_01v8__eta0_diff_30 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_31 = {sky130_fd_pr__pfet_01v8__eta0_diff_31 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_32 = {sky130_fd_pr__pfet_01v8__eta0_diff_32 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_33 = {sky130_fd_pr__pfet_01v8__eta0_diff_33 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_34 = {sky130_fd_pr__pfet_01v8__eta0_diff_34 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_35 = {sky130_fd_pr__pfet_01v8__eta0_diff_35 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_36 = {sky130_fd_pr__pfet_01v8__eta0_diff_36 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_37 = {sky130_fd_pr__pfet_01v8__eta0_diff_37 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_38 = {sky130_fd_pr__pfet_01v8__eta0_diff_38 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_39 = {sky130_fd_pr__pfet_01v8__eta0_diff_39 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_4 = {sky130_fd_pr__pfet_01v8__eta0_diff_4 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_40 = {sky130_fd_pr__pfet_01v8__eta0_diff_40 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_41 = {sky130_fd_pr__pfet_01v8__eta0_diff_41 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_42 = {sky130_fd_pr__pfet_01v8__eta0_diff_42 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_43 = {sky130_fd_pr__pfet_01v8__eta0_diff_43 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_44 = {sky130_fd_pr__pfet_01v8__eta0_diff_44 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_45 = {sky130_fd_pr__pfet_01v8__eta0_diff_45 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_46 = {sky130_fd_pr__pfet_01v8__eta0_diff_46 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_47 = {sky130_fd_pr__pfet_01v8__eta0_diff_47 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_48 = {sky130_fd_pr__pfet_01v8__eta0_diff_48 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_49 = {sky130_fd_pr__pfet_01v8__eta0_diff_49 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_5 = {sky130_fd_pr__pfet_01v8__eta0_diff_5 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_50 = {sky130_fd_pr__pfet_01v8__eta0_diff_50 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_51 = {sky130_fd_pr__pfet_01v8__eta0_diff_51 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_6 = {sky130_fd_pr__pfet_01v8__eta0_diff_6 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_7 = {sky130_fd_pr__pfet_01v8__eta0_diff_7 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_8 = {sky130_fd_pr__pfet_01v8__eta0_diff_8 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__eta0_diff_9 = {sky130_fd_pr__pfet_01v8__eta0_diff_9 + k_pfet_eta0_diff_cd*X_cd + k_pfet_eta0_diff_damage*X_damage + k_pfet_eta0_diff_eot*X_eot + k_pfet_eta0_diff_act*X_act + k_pfet_eta0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_0 = {sky130_fd_pr__pfet_01v8__k2_diff_0 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_1 = {sky130_fd_pr__pfet_01v8__k2_diff_1 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_10 = {sky130_fd_pr__pfet_01v8__k2_diff_10 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_11 = {sky130_fd_pr__pfet_01v8__k2_diff_11 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_12 = {sky130_fd_pr__pfet_01v8__k2_diff_12 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_13 = {sky130_fd_pr__pfet_01v8__k2_diff_13 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_14 = {sky130_fd_pr__pfet_01v8__k2_diff_14 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_15 = {sky130_fd_pr__pfet_01v8__k2_diff_15 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_16 = {sky130_fd_pr__pfet_01v8__k2_diff_16 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_17 = {sky130_fd_pr__pfet_01v8__k2_diff_17 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_18 = {sky130_fd_pr__pfet_01v8__k2_diff_18 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_19 = {sky130_fd_pr__pfet_01v8__k2_diff_19 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_2 = {sky130_fd_pr__pfet_01v8__k2_diff_2 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_20 = {sky130_fd_pr__pfet_01v8__k2_diff_20 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_21 = {sky130_fd_pr__pfet_01v8__k2_diff_21 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_22 = {sky130_fd_pr__pfet_01v8__k2_diff_22 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_23 = {sky130_fd_pr__pfet_01v8__k2_diff_23 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_24 = {sky130_fd_pr__pfet_01v8__k2_diff_24 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_25 = {sky130_fd_pr__pfet_01v8__k2_diff_25 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_26 = {sky130_fd_pr__pfet_01v8__k2_diff_26 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_27 = {sky130_fd_pr__pfet_01v8__k2_diff_27 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_28 = {sky130_fd_pr__pfet_01v8__k2_diff_28 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_29 = {sky130_fd_pr__pfet_01v8__k2_diff_29 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_3 = {sky130_fd_pr__pfet_01v8__k2_diff_3 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_30 = {sky130_fd_pr__pfet_01v8__k2_diff_30 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_31 = {sky130_fd_pr__pfet_01v8__k2_diff_31 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_32 = {sky130_fd_pr__pfet_01v8__k2_diff_32 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_33 = {sky130_fd_pr__pfet_01v8__k2_diff_33 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_34 = {sky130_fd_pr__pfet_01v8__k2_diff_34 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_35 = {sky130_fd_pr__pfet_01v8__k2_diff_35 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_36 = {sky130_fd_pr__pfet_01v8__k2_diff_36 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_37 = {sky130_fd_pr__pfet_01v8__k2_diff_37 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_38 = {sky130_fd_pr__pfet_01v8__k2_diff_38 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_39 = {sky130_fd_pr__pfet_01v8__k2_diff_39 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_4 = {sky130_fd_pr__pfet_01v8__k2_diff_4 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_40 = {sky130_fd_pr__pfet_01v8__k2_diff_40 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_41 = {sky130_fd_pr__pfet_01v8__k2_diff_41 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_42 = {sky130_fd_pr__pfet_01v8__k2_diff_42 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_43 = {sky130_fd_pr__pfet_01v8__k2_diff_43 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_44 = {sky130_fd_pr__pfet_01v8__k2_diff_44 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_45 = {sky130_fd_pr__pfet_01v8__k2_diff_45 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_46 = {sky130_fd_pr__pfet_01v8__k2_diff_46 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_47 = {sky130_fd_pr__pfet_01v8__k2_diff_47 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_48 = {sky130_fd_pr__pfet_01v8__k2_diff_48 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_49 = {sky130_fd_pr__pfet_01v8__k2_diff_49 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_5 = {sky130_fd_pr__pfet_01v8__k2_diff_5 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_50 = {sky130_fd_pr__pfet_01v8__k2_diff_50 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_51 = {sky130_fd_pr__pfet_01v8__k2_diff_51 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_6 = {sky130_fd_pr__pfet_01v8__k2_diff_6 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_7 = {sky130_fd_pr__pfet_01v8__k2_diff_7 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_8 = {sky130_fd_pr__pfet_01v8__k2_diff_8 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__k2_diff_9 = {sky130_fd_pr__pfet_01v8__k2_diff_9 + k_pfet_k2_diff_cd*X_cd + k_pfet_k2_diff_damage*X_damage + k_pfet_k2_diff_eot*X_eot + k_pfet_k2_diff_act*X_act + k_pfet_k2_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_0 = {sky130_fd_pr__pfet_01v8__keta_diff_0 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_1 = {sky130_fd_pr__pfet_01v8__keta_diff_1 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_10 = {sky130_fd_pr__pfet_01v8__keta_diff_10 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_11 = {sky130_fd_pr__pfet_01v8__keta_diff_11 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_12 = {sky130_fd_pr__pfet_01v8__keta_diff_12 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_13 = {sky130_fd_pr__pfet_01v8__keta_diff_13 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_14 = {sky130_fd_pr__pfet_01v8__keta_diff_14 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_15 = {sky130_fd_pr__pfet_01v8__keta_diff_15 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_16 = {sky130_fd_pr__pfet_01v8__keta_diff_16 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_17 = {sky130_fd_pr__pfet_01v8__keta_diff_17 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_18 = {sky130_fd_pr__pfet_01v8__keta_diff_18 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_19 = {sky130_fd_pr__pfet_01v8__keta_diff_19 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_2 = {sky130_fd_pr__pfet_01v8__keta_diff_2 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_20 = {sky130_fd_pr__pfet_01v8__keta_diff_20 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_21 = {sky130_fd_pr__pfet_01v8__keta_diff_21 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_22 = {sky130_fd_pr__pfet_01v8__keta_diff_22 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_23 = {sky130_fd_pr__pfet_01v8__keta_diff_23 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_24 = {sky130_fd_pr__pfet_01v8__keta_diff_24 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_25 = {sky130_fd_pr__pfet_01v8__keta_diff_25 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_26 = {sky130_fd_pr__pfet_01v8__keta_diff_26 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_27 = {sky130_fd_pr__pfet_01v8__keta_diff_27 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_28 = {sky130_fd_pr__pfet_01v8__keta_diff_28 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_29 = {sky130_fd_pr__pfet_01v8__keta_diff_29 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_3 = {sky130_fd_pr__pfet_01v8__keta_diff_3 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_30 = {sky130_fd_pr__pfet_01v8__keta_diff_30 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_31 = {sky130_fd_pr__pfet_01v8__keta_diff_31 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_32 = {sky130_fd_pr__pfet_01v8__keta_diff_32 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_33 = {sky130_fd_pr__pfet_01v8__keta_diff_33 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_34 = {sky130_fd_pr__pfet_01v8__keta_diff_34 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_35 = {sky130_fd_pr__pfet_01v8__keta_diff_35 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_36 = {sky130_fd_pr__pfet_01v8__keta_diff_36 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_37 = {sky130_fd_pr__pfet_01v8__keta_diff_37 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_38 = {sky130_fd_pr__pfet_01v8__keta_diff_38 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_39 = {sky130_fd_pr__pfet_01v8__keta_diff_39 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_4 = {sky130_fd_pr__pfet_01v8__keta_diff_4 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_40 = {sky130_fd_pr__pfet_01v8__keta_diff_40 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_41 = {sky130_fd_pr__pfet_01v8__keta_diff_41 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_42 = {sky130_fd_pr__pfet_01v8__keta_diff_42 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_43 = {sky130_fd_pr__pfet_01v8__keta_diff_43 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_44 = {sky130_fd_pr__pfet_01v8__keta_diff_44 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_45 = {sky130_fd_pr__pfet_01v8__keta_diff_45 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_46 = {sky130_fd_pr__pfet_01v8__keta_diff_46 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_47 = {sky130_fd_pr__pfet_01v8__keta_diff_47 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_48 = {sky130_fd_pr__pfet_01v8__keta_diff_48 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_49 = {sky130_fd_pr__pfet_01v8__keta_diff_49 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_5 = {sky130_fd_pr__pfet_01v8__keta_diff_5 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_50 = {sky130_fd_pr__pfet_01v8__keta_diff_50 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_51 = {sky130_fd_pr__pfet_01v8__keta_diff_51 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_6 = {sky130_fd_pr__pfet_01v8__keta_diff_6 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_7 = {sky130_fd_pr__pfet_01v8__keta_diff_7 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_8 = {sky130_fd_pr__pfet_01v8__keta_diff_8 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__keta_diff_9 = {sky130_fd_pr__pfet_01v8__keta_diff_9 + k_pfet_keta_diff_cd*X_cd + k_pfet_keta_diff_damage*X_damage + k_pfet_keta_diff_eot*X_eot + k_pfet_keta_diff_act*X_act + k_pfet_keta_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_0 = {sky130_fd_pr__pfet_01v8__kt1_diff_0 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_1 = {sky130_fd_pr__pfet_01v8__kt1_diff_1 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_10 = {sky130_fd_pr__pfet_01v8__kt1_diff_10 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_11 = {sky130_fd_pr__pfet_01v8__kt1_diff_11 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_12 = {sky130_fd_pr__pfet_01v8__kt1_diff_12 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_13 = {sky130_fd_pr__pfet_01v8__kt1_diff_13 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_14 = {sky130_fd_pr__pfet_01v8__kt1_diff_14 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_15 = {sky130_fd_pr__pfet_01v8__kt1_diff_15 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_16 = {sky130_fd_pr__pfet_01v8__kt1_diff_16 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_17 = {sky130_fd_pr__pfet_01v8__kt1_diff_17 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_18 = {sky130_fd_pr__pfet_01v8__kt1_diff_18 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_19 = {sky130_fd_pr__pfet_01v8__kt1_diff_19 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_2 = {sky130_fd_pr__pfet_01v8__kt1_diff_2 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_20 = {sky130_fd_pr__pfet_01v8__kt1_diff_20 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_21 = {sky130_fd_pr__pfet_01v8__kt1_diff_21 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_22 = {sky130_fd_pr__pfet_01v8__kt1_diff_22 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_23 = {sky130_fd_pr__pfet_01v8__kt1_diff_23 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_24 = {sky130_fd_pr__pfet_01v8__kt1_diff_24 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_25 = {sky130_fd_pr__pfet_01v8__kt1_diff_25 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_26 = {sky130_fd_pr__pfet_01v8__kt1_diff_26 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_27 = {sky130_fd_pr__pfet_01v8__kt1_diff_27 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_28 = {sky130_fd_pr__pfet_01v8__kt1_diff_28 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_29 = {sky130_fd_pr__pfet_01v8__kt1_diff_29 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_3 = {sky130_fd_pr__pfet_01v8__kt1_diff_3 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_30 = {sky130_fd_pr__pfet_01v8__kt1_diff_30 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_31 = {sky130_fd_pr__pfet_01v8__kt1_diff_31 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_32 = {sky130_fd_pr__pfet_01v8__kt1_diff_32 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_33 = {sky130_fd_pr__pfet_01v8__kt1_diff_33 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_34 = {sky130_fd_pr__pfet_01v8__kt1_diff_34 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_35 = {sky130_fd_pr__pfet_01v8__kt1_diff_35 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_36 = {sky130_fd_pr__pfet_01v8__kt1_diff_36 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_37 = {sky130_fd_pr__pfet_01v8__kt1_diff_37 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_38 = {sky130_fd_pr__pfet_01v8__kt1_diff_38 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_39 = {sky130_fd_pr__pfet_01v8__kt1_diff_39 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_4 = {sky130_fd_pr__pfet_01v8__kt1_diff_4 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_40 = {sky130_fd_pr__pfet_01v8__kt1_diff_40 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_41 = {sky130_fd_pr__pfet_01v8__kt1_diff_41 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_42 = {sky130_fd_pr__pfet_01v8__kt1_diff_42 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_43 = {sky130_fd_pr__pfet_01v8__kt1_diff_43 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_44 = {sky130_fd_pr__pfet_01v8__kt1_diff_44 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_45 = {sky130_fd_pr__pfet_01v8__kt1_diff_45 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_46 = {sky130_fd_pr__pfet_01v8__kt1_diff_46 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_47 = {sky130_fd_pr__pfet_01v8__kt1_diff_47 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_48 = {sky130_fd_pr__pfet_01v8__kt1_diff_48 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_49 = {sky130_fd_pr__pfet_01v8__kt1_diff_49 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_5 = {sky130_fd_pr__pfet_01v8__kt1_diff_5 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_50 = {sky130_fd_pr__pfet_01v8__kt1_diff_50 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_51 = {sky130_fd_pr__pfet_01v8__kt1_diff_51 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_6 = {sky130_fd_pr__pfet_01v8__kt1_diff_6 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_7 = {sky130_fd_pr__pfet_01v8__kt1_diff_7 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_8 = {sky130_fd_pr__pfet_01v8__kt1_diff_8 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__kt1_diff_9 = {sky130_fd_pr__pfet_01v8__kt1_diff_9 + k_pfet_kt1_diff_cd*X_cd + k_pfet_kt1_diff_damage*X_damage + k_pfet_kt1_diff_eot*X_eot + k_pfet_kt1_diff_act*X_act + k_pfet_kt1_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_0 = {sky130_fd_pr__pfet_01v8__nfactor_diff_0 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_1 = {sky130_fd_pr__pfet_01v8__nfactor_diff_1 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_10 = {sky130_fd_pr__pfet_01v8__nfactor_diff_10 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_11 = {sky130_fd_pr__pfet_01v8__nfactor_diff_11 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_12 = {sky130_fd_pr__pfet_01v8__nfactor_diff_12 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_13 = {sky130_fd_pr__pfet_01v8__nfactor_diff_13 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_14 = {sky130_fd_pr__pfet_01v8__nfactor_diff_14 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_15 = {sky130_fd_pr__pfet_01v8__nfactor_diff_15 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_16 = {sky130_fd_pr__pfet_01v8__nfactor_diff_16 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_17 = {sky130_fd_pr__pfet_01v8__nfactor_diff_17 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_18 = {sky130_fd_pr__pfet_01v8__nfactor_diff_18 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_19 = {sky130_fd_pr__pfet_01v8__nfactor_diff_19 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_2 = {sky130_fd_pr__pfet_01v8__nfactor_diff_2 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_20 = {sky130_fd_pr__pfet_01v8__nfactor_diff_20 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_21 = {sky130_fd_pr__pfet_01v8__nfactor_diff_21 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_22 = {sky130_fd_pr__pfet_01v8__nfactor_diff_22 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_23 = {sky130_fd_pr__pfet_01v8__nfactor_diff_23 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_24 = {sky130_fd_pr__pfet_01v8__nfactor_diff_24 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_25 = {sky130_fd_pr__pfet_01v8__nfactor_diff_25 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_26 = {sky130_fd_pr__pfet_01v8__nfactor_diff_26 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_27 = {sky130_fd_pr__pfet_01v8__nfactor_diff_27 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_28 = {sky130_fd_pr__pfet_01v8__nfactor_diff_28 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_29 = {sky130_fd_pr__pfet_01v8__nfactor_diff_29 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_3 = {sky130_fd_pr__pfet_01v8__nfactor_diff_3 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_30 = {sky130_fd_pr__pfet_01v8__nfactor_diff_30 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_31 = {sky130_fd_pr__pfet_01v8__nfactor_diff_31 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_32 = {sky130_fd_pr__pfet_01v8__nfactor_diff_32 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_33 = {sky130_fd_pr__pfet_01v8__nfactor_diff_33 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_34 = {sky130_fd_pr__pfet_01v8__nfactor_diff_34 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_35 = {sky130_fd_pr__pfet_01v8__nfactor_diff_35 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_36 = {sky130_fd_pr__pfet_01v8__nfactor_diff_36 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_37 = {sky130_fd_pr__pfet_01v8__nfactor_diff_37 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_38 = {sky130_fd_pr__pfet_01v8__nfactor_diff_38 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_39 = {sky130_fd_pr__pfet_01v8__nfactor_diff_39 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_4 = {sky130_fd_pr__pfet_01v8__nfactor_diff_4 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_40 = {sky130_fd_pr__pfet_01v8__nfactor_diff_40 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_41 = {sky130_fd_pr__pfet_01v8__nfactor_diff_41 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_42 = {sky130_fd_pr__pfet_01v8__nfactor_diff_42 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_43 = {sky130_fd_pr__pfet_01v8__nfactor_diff_43 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_44 = {sky130_fd_pr__pfet_01v8__nfactor_diff_44 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_45 = {sky130_fd_pr__pfet_01v8__nfactor_diff_45 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_46 = {sky130_fd_pr__pfet_01v8__nfactor_diff_46 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_47 = {sky130_fd_pr__pfet_01v8__nfactor_diff_47 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_48 = {sky130_fd_pr__pfet_01v8__nfactor_diff_48 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_49 = {sky130_fd_pr__pfet_01v8__nfactor_diff_49 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_5 = {sky130_fd_pr__pfet_01v8__nfactor_diff_5 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_50 = {sky130_fd_pr__pfet_01v8__nfactor_diff_50 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_51 = {sky130_fd_pr__pfet_01v8__nfactor_diff_51 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_6 = {sky130_fd_pr__pfet_01v8__nfactor_diff_6 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_7 = {sky130_fd_pr__pfet_01v8__nfactor_diff_7 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_8 = {sky130_fd_pr__pfet_01v8__nfactor_diff_8 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__nfactor_diff_9 = {sky130_fd_pr__pfet_01v8__nfactor_diff_9 + k_pfet_nfactor_diff_cd*X_cd + k_pfet_nfactor_diff_damage*X_damage + k_pfet_nfactor_diff_eot*X_eot + k_pfet_nfactor_diff_act*X_act + k_pfet_nfactor_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_0 = {sky130_fd_pr__pfet_01v8__pclm_diff_0 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_1 = {sky130_fd_pr__pfet_01v8__pclm_diff_1 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_10 = {sky130_fd_pr__pfet_01v8__pclm_diff_10 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_11 = {sky130_fd_pr__pfet_01v8__pclm_diff_11 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_12 = {sky130_fd_pr__pfet_01v8__pclm_diff_12 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_13 = {sky130_fd_pr__pfet_01v8__pclm_diff_13 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_14 = {sky130_fd_pr__pfet_01v8__pclm_diff_14 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_15 = {sky130_fd_pr__pfet_01v8__pclm_diff_15 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_16 = {sky130_fd_pr__pfet_01v8__pclm_diff_16 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_17 = {sky130_fd_pr__pfet_01v8__pclm_diff_17 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_18 = {sky130_fd_pr__pfet_01v8__pclm_diff_18 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_19 = {sky130_fd_pr__pfet_01v8__pclm_diff_19 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_2 = {sky130_fd_pr__pfet_01v8__pclm_diff_2 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_20 = {sky130_fd_pr__pfet_01v8__pclm_diff_20 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_21 = {sky130_fd_pr__pfet_01v8__pclm_diff_21 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_22 = {sky130_fd_pr__pfet_01v8__pclm_diff_22 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_23 = {sky130_fd_pr__pfet_01v8__pclm_diff_23 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_24 = {sky130_fd_pr__pfet_01v8__pclm_diff_24 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_25 = {sky130_fd_pr__pfet_01v8__pclm_diff_25 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_26 = {sky130_fd_pr__pfet_01v8__pclm_diff_26 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_27 = {sky130_fd_pr__pfet_01v8__pclm_diff_27 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_28 = {sky130_fd_pr__pfet_01v8__pclm_diff_28 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_29 = {sky130_fd_pr__pfet_01v8__pclm_diff_29 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_3 = {sky130_fd_pr__pfet_01v8__pclm_diff_3 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_30 = {sky130_fd_pr__pfet_01v8__pclm_diff_30 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_31 = {sky130_fd_pr__pfet_01v8__pclm_diff_31 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_32 = {sky130_fd_pr__pfet_01v8__pclm_diff_32 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_33 = {sky130_fd_pr__pfet_01v8__pclm_diff_33 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_34 = {sky130_fd_pr__pfet_01v8__pclm_diff_34 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_35 = {sky130_fd_pr__pfet_01v8__pclm_diff_35 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_36 = {sky130_fd_pr__pfet_01v8__pclm_diff_36 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_37 = {sky130_fd_pr__pfet_01v8__pclm_diff_37 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_38 = {sky130_fd_pr__pfet_01v8__pclm_diff_38 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_39 = {sky130_fd_pr__pfet_01v8__pclm_diff_39 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_4 = {sky130_fd_pr__pfet_01v8__pclm_diff_4 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_40 = {sky130_fd_pr__pfet_01v8__pclm_diff_40 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_41 = {sky130_fd_pr__pfet_01v8__pclm_diff_41 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_42 = {sky130_fd_pr__pfet_01v8__pclm_diff_42 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_43 = {sky130_fd_pr__pfet_01v8__pclm_diff_43 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_44 = {sky130_fd_pr__pfet_01v8__pclm_diff_44 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_45 = {sky130_fd_pr__pfet_01v8__pclm_diff_45 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_46 = {sky130_fd_pr__pfet_01v8__pclm_diff_46 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_47 = {sky130_fd_pr__pfet_01v8__pclm_diff_47 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_48 = {sky130_fd_pr__pfet_01v8__pclm_diff_48 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_49 = {sky130_fd_pr__pfet_01v8__pclm_diff_49 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_5 = {sky130_fd_pr__pfet_01v8__pclm_diff_5 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_50 = {sky130_fd_pr__pfet_01v8__pclm_diff_50 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_51 = {sky130_fd_pr__pfet_01v8__pclm_diff_51 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_6 = {sky130_fd_pr__pfet_01v8__pclm_diff_6 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_7 = {sky130_fd_pr__pfet_01v8__pclm_diff_7 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_8 = {sky130_fd_pr__pfet_01v8__pclm_diff_8 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pclm_diff_9 = {sky130_fd_pr__pfet_01v8__pclm_diff_9 + k_pfet_pclm_diff_cd*X_cd + k_pfet_pclm_diff_damage*X_damage + k_pfet_pclm_diff_eot*X_eot + k_pfet_pclm_diff_act*X_act + k_pfet_pclm_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_0 = {sky130_fd_pr__pfet_01v8__pdits_diff_0 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_1 = {sky130_fd_pr__pfet_01v8__pdits_diff_1 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_10 = {sky130_fd_pr__pfet_01v8__pdits_diff_10 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_11 = {sky130_fd_pr__pfet_01v8__pdits_diff_11 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_12 = {sky130_fd_pr__pfet_01v8__pdits_diff_12 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_13 = {sky130_fd_pr__pfet_01v8__pdits_diff_13 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_14 = {sky130_fd_pr__pfet_01v8__pdits_diff_14 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_15 = {sky130_fd_pr__pfet_01v8__pdits_diff_15 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_16 = {sky130_fd_pr__pfet_01v8__pdits_diff_16 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_17 = {sky130_fd_pr__pfet_01v8__pdits_diff_17 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_18 = {sky130_fd_pr__pfet_01v8__pdits_diff_18 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_19 = {sky130_fd_pr__pfet_01v8__pdits_diff_19 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_2 = {sky130_fd_pr__pfet_01v8__pdits_diff_2 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_20 = {sky130_fd_pr__pfet_01v8__pdits_diff_20 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_21 = {sky130_fd_pr__pfet_01v8__pdits_diff_21 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_22 = {sky130_fd_pr__pfet_01v8__pdits_diff_22 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_23 = {sky130_fd_pr__pfet_01v8__pdits_diff_23 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_24 = {sky130_fd_pr__pfet_01v8__pdits_diff_24 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_25 = {sky130_fd_pr__pfet_01v8__pdits_diff_25 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_26 = {sky130_fd_pr__pfet_01v8__pdits_diff_26 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_27 = {sky130_fd_pr__pfet_01v8__pdits_diff_27 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_28 = {sky130_fd_pr__pfet_01v8__pdits_diff_28 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_29 = {sky130_fd_pr__pfet_01v8__pdits_diff_29 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_3 = {sky130_fd_pr__pfet_01v8__pdits_diff_3 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_30 = {sky130_fd_pr__pfet_01v8__pdits_diff_30 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_31 = {sky130_fd_pr__pfet_01v8__pdits_diff_31 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_32 = {sky130_fd_pr__pfet_01v8__pdits_diff_32 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_33 = {sky130_fd_pr__pfet_01v8__pdits_diff_33 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_34 = {sky130_fd_pr__pfet_01v8__pdits_diff_34 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_35 = {sky130_fd_pr__pfet_01v8__pdits_diff_35 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_36 = {sky130_fd_pr__pfet_01v8__pdits_diff_36 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_37 = {sky130_fd_pr__pfet_01v8__pdits_diff_37 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_38 = {sky130_fd_pr__pfet_01v8__pdits_diff_38 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_39 = {sky130_fd_pr__pfet_01v8__pdits_diff_39 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_4 = {sky130_fd_pr__pfet_01v8__pdits_diff_4 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_40 = {sky130_fd_pr__pfet_01v8__pdits_diff_40 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_41 = {sky130_fd_pr__pfet_01v8__pdits_diff_41 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_42 = {sky130_fd_pr__pfet_01v8__pdits_diff_42 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_43 = {sky130_fd_pr__pfet_01v8__pdits_diff_43 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_44 = {sky130_fd_pr__pfet_01v8__pdits_diff_44 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_45 = {sky130_fd_pr__pfet_01v8__pdits_diff_45 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_46 = {sky130_fd_pr__pfet_01v8__pdits_diff_46 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_47 = {sky130_fd_pr__pfet_01v8__pdits_diff_47 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_48 = {sky130_fd_pr__pfet_01v8__pdits_diff_48 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_49 = {sky130_fd_pr__pfet_01v8__pdits_diff_49 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_5 = {sky130_fd_pr__pfet_01v8__pdits_diff_5 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_50 = {sky130_fd_pr__pfet_01v8__pdits_diff_50 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_51 = {sky130_fd_pr__pfet_01v8__pdits_diff_51 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_6 = {sky130_fd_pr__pfet_01v8__pdits_diff_6 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_7 = {sky130_fd_pr__pfet_01v8__pdits_diff_7 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_8 = {sky130_fd_pr__pfet_01v8__pdits_diff_8 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pdits_diff_9 = {sky130_fd_pr__pfet_01v8__pdits_diff_9 + k_pfet_pdits_diff_cd*X_cd + k_pfet_pdits_diff_damage*X_damage + k_pfet_pdits_diff_eot*X_eot + k_pfet_pdits_diff_act*X_act + k_pfet_pdits_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_0 = {sky130_fd_pr__pfet_01v8__pditsd_diff_0 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_1 = {sky130_fd_pr__pfet_01v8__pditsd_diff_1 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_10 = {sky130_fd_pr__pfet_01v8__pditsd_diff_10 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_11 = {sky130_fd_pr__pfet_01v8__pditsd_diff_11 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_12 = {sky130_fd_pr__pfet_01v8__pditsd_diff_12 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_13 = {sky130_fd_pr__pfet_01v8__pditsd_diff_13 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_14 = {sky130_fd_pr__pfet_01v8__pditsd_diff_14 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_15 = {sky130_fd_pr__pfet_01v8__pditsd_diff_15 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_16 = {sky130_fd_pr__pfet_01v8__pditsd_diff_16 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_17 = {sky130_fd_pr__pfet_01v8__pditsd_diff_17 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_18 = {sky130_fd_pr__pfet_01v8__pditsd_diff_18 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_19 = {sky130_fd_pr__pfet_01v8__pditsd_diff_19 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_2 = {sky130_fd_pr__pfet_01v8__pditsd_diff_2 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_20 = {sky130_fd_pr__pfet_01v8__pditsd_diff_20 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_21 = {sky130_fd_pr__pfet_01v8__pditsd_diff_21 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_22 = {sky130_fd_pr__pfet_01v8__pditsd_diff_22 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_23 = {sky130_fd_pr__pfet_01v8__pditsd_diff_23 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_24 = {sky130_fd_pr__pfet_01v8__pditsd_diff_24 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_25 = {sky130_fd_pr__pfet_01v8__pditsd_diff_25 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_26 = {sky130_fd_pr__pfet_01v8__pditsd_diff_26 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_27 = {sky130_fd_pr__pfet_01v8__pditsd_diff_27 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_28 = {sky130_fd_pr__pfet_01v8__pditsd_diff_28 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_29 = {sky130_fd_pr__pfet_01v8__pditsd_diff_29 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_3 = {sky130_fd_pr__pfet_01v8__pditsd_diff_3 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_30 = {sky130_fd_pr__pfet_01v8__pditsd_diff_30 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_31 = {sky130_fd_pr__pfet_01v8__pditsd_diff_31 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_32 = {sky130_fd_pr__pfet_01v8__pditsd_diff_32 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_33 = {sky130_fd_pr__pfet_01v8__pditsd_diff_33 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_34 = {sky130_fd_pr__pfet_01v8__pditsd_diff_34 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_35 = {sky130_fd_pr__pfet_01v8__pditsd_diff_35 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_36 = {sky130_fd_pr__pfet_01v8__pditsd_diff_36 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_37 = {sky130_fd_pr__pfet_01v8__pditsd_diff_37 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_38 = {sky130_fd_pr__pfet_01v8__pditsd_diff_38 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_39 = {sky130_fd_pr__pfet_01v8__pditsd_diff_39 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_4 = {sky130_fd_pr__pfet_01v8__pditsd_diff_4 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_40 = {sky130_fd_pr__pfet_01v8__pditsd_diff_40 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_41 = {sky130_fd_pr__pfet_01v8__pditsd_diff_41 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_42 = {sky130_fd_pr__pfet_01v8__pditsd_diff_42 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_43 = {sky130_fd_pr__pfet_01v8__pditsd_diff_43 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_44 = {sky130_fd_pr__pfet_01v8__pditsd_diff_44 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_45 = {sky130_fd_pr__pfet_01v8__pditsd_diff_45 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_46 = {sky130_fd_pr__pfet_01v8__pditsd_diff_46 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_47 = {sky130_fd_pr__pfet_01v8__pditsd_diff_47 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_48 = {sky130_fd_pr__pfet_01v8__pditsd_diff_48 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_49 = {sky130_fd_pr__pfet_01v8__pditsd_diff_49 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_5 = {sky130_fd_pr__pfet_01v8__pditsd_diff_5 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_50 = {sky130_fd_pr__pfet_01v8__pditsd_diff_50 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_51 = {sky130_fd_pr__pfet_01v8__pditsd_diff_51 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_6 = {sky130_fd_pr__pfet_01v8__pditsd_diff_6 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_7 = {sky130_fd_pr__pfet_01v8__pditsd_diff_7 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_8 = {sky130_fd_pr__pfet_01v8__pditsd_diff_8 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__pditsd_diff_9 = {sky130_fd_pr__pfet_01v8__pditsd_diff_9 + k_pfet_pditsd_diff_cd*X_cd + k_pfet_pditsd_diff_damage*X_damage + k_pfet_pditsd_diff_eot*X_eot + k_pfet_pditsd_diff_act*X_act + k_pfet_pditsd_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_0 = {sky130_fd_pr__pfet_01v8__rdsw_diff_0 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_1 = {sky130_fd_pr__pfet_01v8__rdsw_diff_1 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_10 = {sky130_fd_pr__pfet_01v8__rdsw_diff_10 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_11 = {sky130_fd_pr__pfet_01v8__rdsw_diff_11 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_12 = {sky130_fd_pr__pfet_01v8__rdsw_diff_12 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_13 = {sky130_fd_pr__pfet_01v8__rdsw_diff_13 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_14 = {sky130_fd_pr__pfet_01v8__rdsw_diff_14 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_15 = {sky130_fd_pr__pfet_01v8__rdsw_diff_15 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_16 = {sky130_fd_pr__pfet_01v8__rdsw_diff_16 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_17 = {sky130_fd_pr__pfet_01v8__rdsw_diff_17 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_18 = {sky130_fd_pr__pfet_01v8__rdsw_diff_18 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_19 = {sky130_fd_pr__pfet_01v8__rdsw_diff_19 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_2 = {sky130_fd_pr__pfet_01v8__rdsw_diff_2 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_20 = {sky130_fd_pr__pfet_01v8__rdsw_diff_20 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_21 = {sky130_fd_pr__pfet_01v8__rdsw_diff_21 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_22 = {sky130_fd_pr__pfet_01v8__rdsw_diff_22 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_23 = {sky130_fd_pr__pfet_01v8__rdsw_diff_23 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_24 = {sky130_fd_pr__pfet_01v8__rdsw_diff_24 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_25 = {sky130_fd_pr__pfet_01v8__rdsw_diff_25 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_26 = {sky130_fd_pr__pfet_01v8__rdsw_diff_26 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_27 = {sky130_fd_pr__pfet_01v8__rdsw_diff_27 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_28 = {sky130_fd_pr__pfet_01v8__rdsw_diff_28 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_29 = {sky130_fd_pr__pfet_01v8__rdsw_diff_29 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_3 = {sky130_fd_pr__pfet_01v8__rdsw_diff_3 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_30 = {sky130_fd_pr__pfet_01v8__rdsw_diff_30 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_31 = {sky130_fd_pr__pfet_01v8__rdsw_diff_31 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_32 = {sky130_fd_pr__pfet_01v8__rdsw_diff_32 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_33 = {sky130_fd_pr__pfet_01v8__rdsw_diff_33 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_34 = {sky130_fd_pr__pfet_01v8__rdsw_diff_34 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_35 = {sky130_fd_pr__pfet_01v8__rdsw_diff_35 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_36 = {sky130_fd_pr__pfet_01v8__rdsw_diff_36 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_37 = {sky130_fd_pr__pfet_01v8__rdsw_diff_37 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_38 = {sky130_fd_pr__pfet_01v8__rdsw_diff_38 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_39 = {sky130_fd_pr__pfet_01v8__rdsw_diff_39 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_4 = {sky130_fd_pr__pfet_01v8__rdsw_diff_4 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_40 = {sky130_fd_pr__pfet_01v8__rdsw_diff_40 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_41 = {sky130_fd_pr__pfet_01v8__rdsw_diff_41 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_42 = {sky130_fd_pr__pfet_01v8__rdsw_diff_42 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_43 = {sky130_fd_pr__pfet_01v8__rdsw_diff_43 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_44 = {sky130_fd_pr__pfet_01v8__rdsw_diff_44 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_45 = {sky130_fd_pr__pfet_01v8__rdsw_diff_45 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_46 = {sky130_fd_pr__pfet_01v8__rdsw_diff_46 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_47 = {sky130_fd_pr__pfet_01v8__rdsw_diff_47 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_48 = {sky130_fd_pr__pfet_01v8__rdsw_diff_48 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_49 = {sky130_fd_pr__pfet_01v8__rdsw_diff_49 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_5 = {sky130_fd_pr__pfet_01v8__rdsw_diff_5 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_50 = {sky130_fd_pr__pfet_01v8__rdsw_diff_50 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_51 = {sky130_fd_pr__pfet_01v8__rdsw_diff_51 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_6 = {sky130_fd_pr__pfet_01v8__rdsw_diff_6 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_7 = {sky130_fd_pr__pfet_01v8__rdsw_diff_7 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_8 = {sky130_fd_pr__pfet_01v8__rdsw_diff_8 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__rdsw_diff_9 = {sky130_fd_pr__pfet_01v8__rdsw_diff_9 + k_pfet_rdsw_diff_cd*X_cd + k_pfet_rdsw_diff_damage*X_damage + k_pfet_rdsw_diff_eot*X_eot + k_pfet_rdsw_diff_act*X_act + k_pfet_rdsw_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_0 = {sky130_fd_pr__pfet_01v8__tvoff_diff_0 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_1 = {sky130_fd_pr__pfet_01v8__tvoff_diff_1 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_10 = {sky130_fd_pr__pfet_01v8__tvoff_diff_10 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_11 = {sky130_fd_pr__pfet_01v8__tvoff_diff_11 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_12 = {sky130_fd_pr__pfet_01v8__tvoff_diff_12 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_13 = {sky130_fd_pr__pfet_01v8__tvoff_diff_13 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_14 = {sky130_fd_pr__pfet_01v8__tvoff_diff_14 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_15 = {sky130_fd_pr__pfet_01v8__tvoff_diff_15 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_16 = {sky130_fd_pr__pfet_01v8__tvoff_diff_16 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_17 = {sky130_fd_pr__pfet_01v8__tvoff_diff_17 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_18 = {sky130_fd_pr__pfet_01v8__tvoff_diff_18 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_19 = {sky130_fd_pr__pfet_01v8__tvoff_diff_19 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_2 = {sky130_fd_pr__pfet_01v8__tvoff_diff_2 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_20 = {sky130_fd_pr__pfet_01v8__tvoff_diff_20 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_21 = {sky130_fd_pr__pfet_01v8__tvoff_diff_21 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_22 = {sky130_fd_pr__pfet_01v8__tvoff_diff_22 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_23 = {sky130_fd_pr__pfet_01v8__tvoff_diff_23 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_24 = {sky130_fd_pr__pfet_01v8__tvoff_diff_24 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_25 = {sky130_fd_pr__pfet_01v8__tvoff_diff_25 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_26 = {sky130_fd_pr__pfet_01v8__tvoff_diff_26 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_27 = {sky130_fd_pr__pfet_01v8__tvoff_diff_27 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_28 = {sky130_fd_pr__pfet_01v8__tvoff_diff_28 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_29 = {sky130_fd_pr__pfet_01v8__tvoff_diff_29 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_3 = {sky130_fd_pr__pfet_01v8__tvoff_diff_3 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_30 = {sky130_fd_pr__pfet_01v8__tvoff_diff_30 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_31 = {sky130_fd_pr__pfet_01v8__tvoff_diff_31 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_32 = {sky130_fd_pr__pfet_01v8__tvoff_diff_32 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_33 = {sky130_fd_pr__pfet_01v8__tvoff_diff_33 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_34 = {sky130_fd_pr__pfet_01v8__tvoff_diff_34 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_35 = {sky130_fd_pr__pfet_01v8__tvoff_diff_35 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_36 = {sky130_fd_pr__pfet_01v8__tvoff_diff_36 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_37 = {sky130_fd_pr__pfet_01v8__tvoff_diff_37 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_38 = {sky130_fd_pr__pfet_01v8__tvoff_diff_38 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_39 = {sky130_fd_pr__pfet_01v8__tvoff_diff_39 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_4 = {sky130_fd_pr__pfet_01v8__tvoff_diff_4 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_40 = {sky130_fd_pr__pfet_01v8__tvoff_diff_40 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_41 = {sky130_fd_pr__pfet_01v8__tvoff_diff_41 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_42 = {sky130_fd_pr__pfet_01v8__tvoff_diff_42 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_43 = {sky130_fd_pr__pfet_01v8__tvoff_diff_43 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_44 = {sky130_fd_pr__pfet_01v8__tvoff_diff_44 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_45 = {sky130_fd_pr__pfet_01v8__tvoff_diff_45 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_46 = {sky130_fd_pr__pfet_01v8__tvoff_diff_46 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_47 = {sky130_fd_pr__pfet_01v8__tvoff_diff_47 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_48 = {sky130_fd_pr__pfet_01v8__tvoff_diff_48 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_49 = {sky130_fd_pr__pfet_01v8__tvoff_diff_49 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_5 = {sky130_fd_pr__pfet_01v8__tvoff_diff_5 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_50 = {sky130_fd_pr__pfet_01v8__tvoff_diff_50 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_51 = {sky130_fd_pr__pfet_01v8__tvoff_diff_51 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_6 = {sky130_fd_pr__pfet_01v8__tvoff_diff_6 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_7 = {sky130_fd_pr__pfet_01v8__tvoff_diff_7 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_8 = {sky130_fd_pr__pfet_01v8__tvoff_diff_8 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__tvoff_diff_9 = {sky130_fd_pr__pfet_01v8__tvoff_diff_9 + k_pfet_tvoff_diff_cd*X_cd + k_pfet_tvoff_diff_damage*X_damage + k_pfet_tvoff_diff_eot*X_eot + k_pfet_tvoff_diff_act*X_act + k_pfet_tvoff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_0 = {sky130_fd_pr__pfet_01v8__u0_diff_0 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_1 = {sky130_fd_pr__pfet_01v8__u0_diff_1 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_10 = {sky130_fd_pr__pfet_01v8__u0_diff_10 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_11 = {sky130_fd_pr__pfet_01v8__u0_diff_11 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_12 = {sky130_fd_pr__pfet_01v8__u0_diff_12 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_13 = {sky130_fd_pr__pfet_01v8__u0_diff_13 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_14 = {sky130_fd_pr__pfet_01v8__u0_diff_14 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_15 = {sky130_fd_pr__pfet_01v8__u0_diff_15 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_16 = {sky130_fd_pr__pfet_01v8__u0_diff_16 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_17 = {sky130_fd_pr__pfet_01v8__u0_diff_17 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_18 = {sky130_fd_pr__pfet_01v8__u0_diff_18 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_19 = {sky130_fd_pr__pfet_01v8__u0_diff_19 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_2 = {sky130_fd_pr__pfet_01v8__u0_diff_2 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_20 = {sky130_fd_pr__pfet_01v8__u0_diff_20 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_21 = {sky130_fd_pr__pfet_01v8__u0_diff_21 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_22 = {sky130_fd_pr__pfet_01v8__u0_diff_22 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_23 = {sky130_fd_pr__pfet_01v8__u0_diff_23 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_24 = {sky130_fd_pr__pfet_01v8__u0_diff_24 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_25 = {sky130_fd_pr__pfet_01v8__u0_diff_25 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_26 = {sky130_fd_pr__pfet_01v8__u0_diff_26 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_27 = {sky130_fd_pr__pfet_01v8__u0_diff_27 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_28 = {sky130_fd_pr__pfet_01v8__u0_diff_28 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_29 = {sky130_fd_pr__pfet_01v8__u0_diff_29 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_3 = {sky130_fd_pr__pfet_01v8__u0_diff_3 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_30 = {sky130_fd_pr__pfet_01v8__u0_diff_30 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_31 = {sky130_fd_pr__pfet_01v8__u0_diff_31 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_32 = {sky130_fd_pr__pfet_01v8__u0_diff_32 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_33 = {sky130_fd_pr__pfet_01v8__u0_diff_33 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_34 = {sky130_fd_pr__pfet_01v8__u0_diff_34 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_35 = {sky130_fd_pr__pfet_01v8__u0_diff_35 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_36 = {sky130_fd_pr__pfet_01v8__u0_diff_36 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_37 = {sky130_fd_pr__pfet_01v8__u0_diff_37 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_38 = {sky130_fd_pr__pfet_01v8__u0_diff_38 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_39 = {sky130_fd_pr__pfet_01v8__u0_diff_39 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_4 = {sky130_fd_pr__pfet_01v8__u0_diff_4 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_40 = {sky130_fd_pr__pfet_01v8__u0_diff_40 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_41 = {sky130_fd_pr__pfet_01v8__u0_diff_41 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_42 = {sky130_fd_pr__pfet_01v8__u0_diff_42 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_43 = {sky130_fd_pr__pfet_01v8__u0_diff_43 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_44 = {sky130_fd_pr__pfet_01v8__u0_diff_44 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_45 = {sky130_fd_pr__pfet_01v8__u0_diff_45 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_46 = {sky130_fd_pr__pfet_01v8__u0_diff_46 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_47 = {sky130_fd_pr__pfet_01v8__u0_diff_47 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_48 = {sky130_fd_pr__pfet_01v8__u0_diff_48 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_49 = {sky130_fd_pr__pfet_01v8__u0_diff_49 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_5 = {sky130_fd_pr__pfet_01v8__u0_diff_5 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_50 = {sky130_fd_pr__pfet_01v8__u0_diff_50 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_51 = {sky130_fd_pr__pfet_01v8__u0_diff_51 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_6 = {sky130_fd_pr__pfet_01v8__u0_diff_6 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_7 = {sky130_fd_pr__pfet_01v8__u0_diff_7 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_8 = {sky130_fd_pr__pfet_01v8__u0_diff_8 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__u0_diff_9 = {sky130_fd_pr__pfet_01v8__u0_diff_9 + k_pfet_u0_diff_cd*X_cd + k_pfet_u0_diff_damage*X_damage + k_pfet_u0_diff_eot*X_eot + k_pfet_u0_diff_act*X_act + k_pfet_u0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_0 = {sky130_fd_pr__pfet_01v8__ua_diff_0 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_1 = {sky130_fd_pr__pfet_01v8__ua_diff_1 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_10 = {sky130_fd_pr__pfet_01v8__ua_diff_10 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_11 = {sky130_fd_pr__pfet_01v8__ua_diff_11 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_12 = {sky130_fd_pr__pfet_01v8__ua_diff_12 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_13 = {sky130_fd_pr__pfet_01v8__ua_diff_13 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_14 = {sky130_fd_pr__pfet_01v8__ua_diff_14 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_15 = {sky130_fd_pr__pfet_01v8__ua_diff_15 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_16 = {sky130_fd_pr__pfet_01v8__ua_diff_16 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_17 = {sky130_fd_pr__pfet_01v8__ua_diff_17 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_18 = {sky130_fd_pr__pfet_01v8__ua_diff_18 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_19 = {sky130_fd_pr__pfet_01v8__ua_diff_19 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_2 = {sky130_fd_pr__pfet_01v8__ua_diff_2 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_20 = {sky130_fd_pr__pfet_01v8__ua_diff_20 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_21 = {sky130_fd_pr__pfet_01v8__ua_diff_21 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_22 = {sky130_fd_pr__pfet_01v8__ua_diff_22 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_23 = {sky130_fd_pr__pfet_01v8__ua_diff_23 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_24 = {sky130_fd_pr__pfet_01v8__ua_diff_24 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_25 = {sky130_fd_pr__pfet_01v8__ua_diff_25 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_26 = {sky130_fd_pr__pfet_01v8__ua_diff_26 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_27 = {sky130_fd_pr__pfet_01v8__ua_diff_27 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_28 = {sky130_fd_pr__pfet_01v8__ua_diff_28 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_29 = {sky130_fd_pr__pfet_01v8__ua_diff_29 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_3 = {sky130_fd_pr__pfet_01v8__ua_diff_3 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_30 = {sky130_fd_pr__pfet_01v8__ua_diff_30 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_31 = {sky130_fd_pr__pfet_01v8__ua_diff_31 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_32 = {sky130_fd_pr__pfet_01v8__ua_diff_32 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_33 = {sky130_fd_pr__pfet_01v8__ua_diff_33 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_34 = {sky130_fd_pr__pfet_01v8__ua_diff_34 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_35 = {sky130_fd_pr__pfet_01v8__ua_diff_35 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_36 = {sky130_fd_pr__pfet_01v8__ua_diff_36 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_37 = {sky130_fd_pr__pfet_01v8__ua_diff_37 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_38 = {sky130_fd_pr__pfet_01v8__ua_diff_38 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_39 = {sky130_fd_pr__pfet_01v8__ua_diff_39 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_4 = {sky130_fd_pr__pfet_01v8__ua_diff_4 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_40 = {sky130_fd_pr__pfet_01v8__ua_diff_40 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_41 = {sky130_fd_pr__pfet_01v8__ua_diff_41 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_42 = {sky130_fd_pr__pfet_01v8__ua_diff_42 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_43 = {sky130_fd_pr__pfet_01v8__ua_diff_43 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_44 = {sky130_fd_pr__pfet_01v8__ua_diff_44 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_45 = {sky130_fd_pr__pfet_01v8__ua_diff_45 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_46 = {sky130_fd_pr__pfet_01v8__ua_diff_46 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_47 = {sky130_fd_pr__pfet_01v8__ua_diff_47 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_48 = {sky130_fd_pr__pfet_01v8__ua_diff_48 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_49 = {sky130_fd_pr__pfet_01v8__ua_diff_49 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_5 = {sky130_fd_pr__pfet_01v8__ua_diff_5 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_50 = {sky130_fd_pr__pfet_01v8__ua_diff_50 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_51 = {sky130_fd_pr__pfet_01v8__ua_diff_51 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_6 = {sky130_fd_pr__pfet_01v8__ua_diff_6 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_7 = {sky130_fd_pr__pfet_01v8__ua_diff_7 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_8 = {sky130_fd_pr__pfet_01v8__ua_diff_8 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ua_diff_9 = {sky130_fd_pr__pfet_01v8__ua_diff_9 + k_pfet_ua_diff_cd*X_cd + k_pfet_ua_diff_damage*X_damage + k_pfet_ua_diff_eot*X_eot + k_pfet_ua_diff_act*X_act + k_pfet_ua_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_0 = {sky130_fd_pr__pfet_01v8__ub_diff_0 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_1 = {sky130_fd_pr__pfet_01v8__ub_diff_1 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_10 = {sky130_fd_pr__pfet_01v8__ub_diff_10 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_11 = {sky130_fd_pr__pfet_01v8__ub_diff_11 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_12 = {sky130_fd_pr__pfet_01v8__ub_diff_12 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_13 = {sky130_fd_pr__pfet_01v8__ub_diff_13 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_14 = {sky130_fd_pr__pfet_01v8__ub_diff_14 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_15 = {sky130_fd_pr__pfet_01v8__ub_diff_15 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_16 = {sky130_fd_pr__pfet_01v8__ub_diff_16 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_17 = {sky130_fd_pr__pfet_01v8__ub_diff_17 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_18 = {sky130_fd_pr__pfet_01v8__ub_diff_18 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_19 = {sky130_fd_pr__pfet_01v8__ub_diff_19 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_2 = {sky130_fd_pr__pfet_01v8__ub_diff_2 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_20 = {sky130_fd_pr__pfet_01v8__ub_diff_20 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_21 = {sky130_fd_pr__pfet_01v8__ub_diff_21 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_22 = {sky130_fd_pr__pfet_01v8__ub_diff_22 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_23 = {sky130_fd_pr__pfet_01v8__ub_diff_23 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_24 = {sky130_fd_pr__pfet_01v8__ub_diff_24 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_25 = {sky130_fd_pr__pfet_01v8__ub_diff_25 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_26 = {sky130_fd_pr__pfet_01v8__ub_diff_26 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_27 = {sky130_fd_pr__pfet_01v8__ub_diff_27 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_28 = {sky130_fd_pr__pfet_01v8__ub_diff_28 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_29 = {sky130_fd_pr__pfet_01v8__ub_diff_29 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_3 = {sky130_fd_pr__pfet_01v8__ub_diff_3 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_30 = {sky130_fd_pr__pfet_01v8__ub_diff_30 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_31 = {sky130_fd_pr__pfet_01v8__ub_diff_31 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_32 = {sky130_fd_pr__pfet_01v8__ub_diff_32 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_33 = {sky130_fd_pr__pfet_01v8__ub_diff_33 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_34 = {sky130_fd_pr__pfet_01v8__ub_diff_34 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_35 = {sky130_fd_pr__pfet_01v8__ub_diff_35 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_36 = {sky130_fd_pr__pfet_01v8__ub_diff_36 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_37 = {sky130_fd_pr__pfet_01v8__ub_diff_37 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_38 = {sky130_fd_pr__pfet_01v8__ub_diff_38 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_39 = {sky130_fd_pr__pfet_01v8__ub_diff_39 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_4 = {sky130_fd_pr__pfet_01v8__ub_diff_4 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_40 = {sky130_fd_pr__pfet_01v8__ub_diff_40 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_41 = {sky130_fd_pr__pfet_01v8__ub_diff_41 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_42 = {sky130_fd_pr__pfet_01v8__ub_diff_42 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_43 = {sky130_fd_pr__pfet_01v8__ub_diff_43 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_44 = {sky130_fd_pr__pfet_01v8__ub_diff_44 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_45 = {sky130_fd_pr__pfet_01v8__ub_diff_45 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_46 = {sky130_fd_pr__pfet_01v8__ub_diff_46 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_47 = {sky130_fd_pr__pfet_01v8__ub_diff_47 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_48 = {sky130_fd_pr__pfet_01v8__ub_diff_48 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_49 = {sky130_fd_pr__pfet_01v8__ub_diff_49 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_5 = {sky130_fd_pr__pfet_01v8__ub_diff_5 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_50 = {sky130_fd_pr__pfet_01v8__ub_diff_50 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_51 = {sky130_fd_pr__pfet_01v8__ub_diff_51 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_6 = {sky130_fd_pr__pfet_01v8__ub_diff_6 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_7 = {sky130_fd_pr__pfet_01v8__ub_diff_7 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_8 = {sky130_fd_pr__pfet_01v8__ub_diff_8 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__ub_diff_9 = {sky130_fd_pr__pfet_01v8__ub_diff_9 + k_pfet_ub_diff_cd*X_cd + k_pfet_ub_diff_damage*X_damage + k_pfet_ub_diff_eot*X_eot + k_pfet_ub_diff_act*X_act + k_pfet_ub_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_0 = {sky130_fd_pr__pfet_01v8__voff_diff_0 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_1 = {sky130_fd_pr__pfet_01v8__voff_diff_1 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_10 = {sky130_fd_pr__pfet_01v8__voff_diff_10 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_11 = {sky130_fd_pr__pfet_01v8__voff_diff_11 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_12 = {sky130_fd_pr__pfet_01v8__voff_diff_12 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_13 = {sky130_fd_pr__pfet_01v8__voff_diff_13 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_14 = {sky130_fd_pr__pfet_01v8__voff_diff_14 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_15 = {sky130_fd_pr__pfet_01v8__voff_diff_15 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_16 = {sky130_fd_pr__pfet_01v8__voff_diff_16 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_17 = {sky130_fd_pr__pfet_01v8__voff_diff_17 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_18 = {sky130_fd_pr__pfet_01v8__voff_diff_18 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_19 = {sky130_fd_pr__pfet_01v8__voff_diff_19 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_2 = {sky130_fd_pr__pfet_01v8__voff_diff_2 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_20 = {sky130_fd_pr__pfet_01v8__voff_diff_20 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_21 = {sky130_fd_pr__pfet_01v8__voff_diff_21 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_22 = {sky130_fd_pr__pfet_01v8__voff_diff_22 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_23 = {sky130_fd_pr__pfet_01v8__voff_diff_23 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_24 = {sky130_fd_pr__pfet_01v8__voff_diff_24 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_25 = {sky130_fd_pr__pfet_01v8__voff_diff_25 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_26 = {sky130_fd_pr__pfet_01v8__voff_diff_26 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_27 = {sky130_fd_pr__pfet_01v8__voff_diff_27 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_28 = {sky130_fd_pr__pfet_01v8__voff_diff_28 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_29 = {sky130_fd_pr__pfet_01v8__voff_diff_29 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_3 = {sky130_fd_pr__pfet_01v8__voff_diff_3 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_30 = {sky130_fd_pr__pfet_01v8__voff_diff_30 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_31 = {sky130_fd_pr__pfet_01v8__voff_diff_31 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_32 = {sky130_fd_pr__pfet_01v8__voff_diff_32 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_33 = {sky130_fd_pr__pfet_01v8__voff_diff_33 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_34 = {sky130_fd_pr__pfet_01v8__voff_diff_34 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_35 = {sky130_fd_pr__pfet_01v8__voff_diff_35 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_36 = {sky130_fd_pr__pfet_01v8__voff_diff_36 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_37 = {sky130_fd_pr__pfet_01v8__voff_diff_37 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_38 = {sky130_fd_pr__pfet_01v8__voff_diff_38 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_39 = {sky130_fd_pr__pfet_01v8__voff_diff_39 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_4 = {sky130_fd_pr__pfet_01v8__voff_diff_4 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_40 = {sky130_fd_pr__pfet_01v8__voff_diff_40 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_41 = {sky130_fd_pr__pfet_01v8__voff_diff_41 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_42 = {sky130_fd_pr__pfet_01v8__voff_diff_42 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_43 = {sky130_fd_pr__pfet_01v8__voff_diff_43 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_44 = {sky130_fd_pr__pfet_01v8__voff_diff_44 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_45 = {sky130_fd_pr__pfet_01v8__voff_diff_45 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_46 = {sky130_fd_pr__pfet_01v8__voff_diff_46 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_47 = {sky130_fd_pr__pfet_01v8__voff_diff_47 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_48 = {sky130_fd_pr__pfet_01v8__voff_diff_48 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_49 = {sky130_fd_pr__pfet_01v8__voff_diff_49 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_5 = {sky130_fd_pr__pfet_01v8__voff_diff_5 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_50 = {sky130_fd_pr__pfet_01v8__voff_diff_50 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_51 = {sky130_fd_pr__pfet_01v8__voff_diff_51 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_6 = {sky130_fd_pr__pfet_01v8__voff_diff_6 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_7 = {sky130_fd_pr__pfet_01v8__voff_diff_7 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_8 = {sky130_fd_pr__pfet_01v8__voff_diff_8 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__voff_diff_9 = {sky130_fd_pr__pfet_01v8__voff_diff_9 + k_pfet_voff_diff_cd*X_cd + k_pfet_voff_diff_damage*X_damage + k_pfet_voff_diff_eot*X_eot + k_pfet_voff_diff_act*X_act + k_pfet_voff_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_0 = {sky130_fd_pr__pfet_01v8__vsat_diff_0 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_1 = {sky130_fd_pr__pfet_01v8__vsat_diff_1 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_10 = {sky130_fd_pr__pfet_01v8__vsat_diff_10 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_11 = {sky130_fd_pr__pfet_01v8__vsat_diff_11 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_12 = {sky130_fd_pr__pfet_01v8__vsat_diff_12 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_13 = {sky130_fd_pr__pfet_01v8__vsat_diff_13 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_14 = {sky130_fd_pr__pfet_01v8__vsat_diff_14 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_15 = {sky130_fd_pr__pfet_01v8__vsat_diff_15 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_16 = {sky130_fd_pr__pfet_01v8__vsat_diff_16 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_17 = {sky130_fd_pr__pfet_01v8__vsat_diff_17 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_18 = {sky130_fd_pr__pfet_01v8__vsat_diff_18 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_19 = {sky130_fd_pr__pfet_01v8__vsat_diff_19 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_2 = {sky130_fd_pr__pfet_01v8__vsat_diff_2 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_20 = {sky130_fd_pr__pfet_01v8__vsat_diff_20 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_21 = {sky130_fd_pr__pfet_01v8__vsat_diff_21 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_22 = {sky130_fd_pr__pfet_01v8__vsat_diff_22 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_23 = {sky130_fd_pr__pfet_01v8__vsat_diff_23 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_24 = {sky130_fd_pr__pfet_01v8__vsat_diff_24 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_25 = {sky130_fd_pr__pfet_01v8__vsat_diff_25 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_26 = {sky130_fd_pr__pfet_01v8__vsat_diff_26 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_27 = {sky130_fd_pr__pfet_01v8__vsat_diff_27 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_28 = {sky130_fd_pr__pfet_01v8__vsat_diff_28 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_29 = {sky130_fd_pr__pfet_01v8__vsat_diff_29 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_3 = {sky130_fd_pr__pfet_01v8__vsat_diff_3 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_30 = {sky130_fd_pr__pfet_01v8__vsat_diff_30 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_31 = {sky130_fd_pr__pfet_01v8__vsat_diff_31 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_32 = {sky130_fd_pr__pfet_01v8__vsat_diff_32 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_33 = {sky130_fd_pr__pfet_01v8__vsat_diff_33 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_34 = {sky130_fd_pr__pfet_01v8__vsat_diff_34 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_35 = {sky130_fd_pr__pfet_01v8__vsat_diff_35 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_36 = {sky130_fd_pr__pfet_01v8__vsat_diff_36 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_37 = {sky130_fd_pr__pfet_01v8__vsat_diff_37 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_38 = {sky130_fd_pr__pfet_01v8__vsat_diff_38 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_39 = {sky130_fd_pr__pfet_01v8__vsat_diff_39 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_4 = {sky130_fd_pr__pfet_01v8__vsat_diff_4 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_40 = {sky130_fd_pr__pfet_01v8__vsat_diff_40 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_41 = {sky130_fd_pr__pfet_01v8__vsat_diff_41 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_42 = {sky130_fd_pr__pfet_01v8__vsat_diff_42 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_43 = {sky130_fd_pr__pfet_01v8__vsat_diff_43 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_44 = {sky130_fd_pr__pfet_01v8__vsat_diff_44 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_45 = {sky130_fd_pr__pfet_01v8__vsat_diff_45 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_46 = {sky130_fd_pr__pfet_01v8__vsat_diff_46 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_47 = {sky130_fd_pr__pfet_01v8__vsat_diff_47 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_48 = {sky130_fd_pr__pfet_01v8__vsat_diff_48 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_49 = {sky130_fd_pr__pfet_01v8__vsat_diff_49 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_5 = {sky130_fd_pr__pfet_01v8__vsat_diff_5 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_50 = {sky130_fd_pr__pfet_01v8__vsat_diff_50 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_51 = {sky130_fd_pr__pfet_01v8__vsat_diff_51 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_6 = {sky130_fd_pr__pfet_01v8__vsat_diff_6 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_7 = {sky130_fd_pr__pfet_01v8__vsat_diff_7 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_8 = {sky130_fd_pr__pfet_01v8__vsat_diff_8 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vsat_diff_9 = {sky130_fd_pr__pfet_01v8__vsat_diff_9 + k_pfet_vsat_diff_cd*X_cd + k_pfet_vsat_diff_damage*X_damage + k_pfet_vsat_diff_eot*X_eot + k_pfet_vsat_diff_act*X_act + k_pfet_vsat_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_0 = {sky130_fd_pr__pfet_01v8__vth0_diff_0 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_1 = {sky130_fd_pr__pfet_01v8__vth0_diff_1 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_10 = {sky130_fd_pr__pfet_01v8__vth0_diff_10 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_11 = {sky130_fd_pr__pfet_01v8__vth0_diff_11 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_12 = {sky130_fd_pr__pfet_01v8__vth0_diff_12 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_13 = {sky130_fd_pr__pfet_01v8__vth0_diff_13 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_14 = {sky130_fd_pr__pfet_01v8__vth0_diff_14 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_15 = {sky130_fd_pr__pfet_01v8__vth0_diff_15 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_16 = {sky130_fd_pr__pfet_01v8__vth0_diff_16 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_17 = {sky130_fd_pr__pfet_01v8__vth0_diff_17 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_18 = {sky130_fd_pr__pfet_01v8__vth0_diff_18 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_19 = {sky130_fd_pr__pfet_01v8__vth0_diff_19 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_2 = {sky130_fd_pr__pfet_01v8__vth0_diff_2 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_20 = {sky130_fd_pr__pfet_01v8__vth0_diff_20 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_21 = {sky130_fd_pr__pfet_01v8__vth0_diff_21 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_22 = {sky130_fd_pr__pfet_01v8__vth0_diff_22 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_23 = {sky130_fd_pr__pfet_01v8__vth0_diff_23 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_24 = {sky130_fd_pr__pfet_01v8__vth0_diff_24 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_25 = {sky130_fd_pr__pfet_01v8__vth0_diff_25 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_26 = {sky130_fd_pr__pfet_01v8__vth0_diff_26 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_27 = {sky130_fd_pr__pfet_01v8__vth0_diff_27 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_28 = {sky130_fd_pr__pfet_01v8__vth0_diff_28 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_29 = {sky130_fd_pr__pfet_01v8__vth0_diff_29 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_3 = {sky130_fd_pr__pfet_01v8__vth0_diff_3 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_30 = {sky130_fd_pr__pfet_01v8__vth0_diff_30 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_31 = {sky130_fd_pr__pfet_01v8__vth0_diff_31 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_32 = {sky130_fd_pr__pfet_01v8__vth0_diff_32 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_33 = {sky130_fd_pr__pfet_01v8__vth0_diff_33 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_34 = {sky130_fd_pr__pfet_01v8__vth0_diff_34 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_35 = {sky130_fd_pr__pfet_01v8__vth0_diff_35 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_36 = {sky130_fd_pr__pfet_01v8__vth0_diff_36 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_37 = {sky130_fd_pr__pfet_01v8__vth0_diff_37 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_38 = {sky130_fd_pr__pfet_01v8__vth0_diff_38 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_39 = {sky130_fd_pr__pfet_01v8__vth0_diff_39 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_4 = {sky130_fd_pr__pfet_01v8__vth0_diff_4 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_40 = {sky130_fd_pr__pfet_01v8__vth0_diff_40 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_41 = {sky130_fd_pr__pfet_01v8__vth0_diff_41 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_42 = {sky130_fd_pr__pfet_01v8__vth0_diff_42 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_43 = {sky130_fd_pr__pfet_01v8__vth0_diff_43 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_44 = {sky130_fd_pr__pfet_01v8__vth0_diff_44 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_45 = {sky130_fd_pr__pfet_01v8__vth0_diff_45 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_46 = {sky130_fd_pr__pfet_01v8__vth0_diff_46 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_47 = {sky130_fd_pr__pfet_01v8__vth0_diff_47 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_48 = {sky130_fd_pr__pfet_01v8__vth0_diff_48 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_49 = {sky130_fd_pr__pfet_01v8__vth0_diff_49 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_5 = {sky130_fd_pr__pfet_01v8__vth0_diff_5 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_50 = {sky130_fd_pr__pfet_01v8__vth0_diff_50 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_51 = {sky130_fd_pr__pfet_01v8__vth0_diff_51 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_6 = {sky130_fd_pr__pfet_01v8__vth0_diff_6 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_7 = {sky130_fd_pr__pfet_01v8__vth0_diff_7 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_8 = {sky130_fd_pr__pfet_01v8__vth0_diff_8 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}
.param sky130_fd_pr__pfet_01v8__vth0_diff_9 = {sky130_fd_pr__pfet_01v8__vth0_diff_9 + k_pfet_vth0_diff_cd*X_cd + k_pfet_vth0_diff_damage*X_damage + k_pfet_vth0_diff_eot*X_eot + k_pfet_vth0_diff_act*X_act + k_pfet_vth0_diff_rc*X_rc}

* ============================================================
* END ROOT-CAUSE OVERRIDES
* === ROOTCAUSE_UI_END ===
* ============================================================
